
module Register_File_WIDTH32_DEPTH5_1 ( clk, reset, read_enable_1, 
        read_enable_2, write_enable, read_index_1, read_index_2, write_index, 
        write_data, read_data_1, read_data_2 );
  input [4:0] read_index_1;
  input [4:0] read_index_2;
  input [4:0] write_index;
  input [31:0] write_data;
  output [31:0] read_data_1;
  output [31:0] read_data_2;
  input clk, reset, read_enable_1, read_enable_2, write_enable;

  tri   [31:0] read_data_1;
  tri   [31:0] read_data_2;

  TBUFX2 \read_data_1_tri[31]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[31]) );
  TBUFX2 \read_data_1_tri[30]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[30]) );
  TBUFX2 \read_data_1_tri[29]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[29]) );
  TBUFX2 \read_data_1_tri[28]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[28]) );
  TBUFX2 \read_data_1_tri[27]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[27]) );
  TBUFX2 \read_data_1_tri[26]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[26]) );
  TBUFX2 \read_data_1_tri[25]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[25]) );
  TBUFX2 \read_data_1_tri[24]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[24]) );
  TBUFX2 \read_data_1_tri[23]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[23]) );
  TBUFX2 \read_data_1_tri[22]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[22]) );
  TBUFX2 \read_data_1_tri[21]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[21]) );
  TBUFX2 \read_data_1_tri[20]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[20]) );
  TBUFX2 \read_data_1_tri[19]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[19]) );
  TBUFX2 \read_data_1_tri[18]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[18]) );
  TBUFX2 \read_data_1_tri[17]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[17]) );
  TBUFX2 \read_data_1_tri[16]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[16]) );
  TBUFX2 \read_data_1_tri[15]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[15]) );
  TBUFX2 \read_data_1_tri[14]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[14]) );
  TBUFX2 \read_data_1_tri[13]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[13]) );
  TBUFX2 \read_data_1_tri[12]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[12]) );
  TBUFX2 \read_data_1_tri[11]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[11]) );
  TBUFX2 \read_data_1_tri[10]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[10]) );
  TBUFX2 \read_data_1_tri[8]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[8]) );
  TBUFX2 \read_data_1_tri[7]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[7]) );
  TBUFX2 \read_data_1_tri[6]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[6]) );
  TBUFX2 \read_data_1_tri[5]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[5]) );
  TBUFX2 \read_data_1_tri[4]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[4]) );
  TBUFX2 \read_data_1_tri[3]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[3]) );
  TBUFX2 \read_data_1_tri[2]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[2]) );
  TBUFX2 \read_data_1_tri[1]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[1]) );
  TBUFX2 \read_data_1_tri[0]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[0]) );
  TBUFX2 \read_data_2_tri[31]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[31]) );
  TBUFX2 \read_data_2_tri[30]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[30]) );
  TBUFX2 \read_data_2_tri[28]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[28]) );
  TBUFX2 \read_data_2_tri[27]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[27]) );
  TBUFX2 \read_data_2_tri[26]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[26]) );
  TBUFX2 \read_data_2_tri[25]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[25]) );
  TBUFX2 \read_data_2_tri[24]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[24]) );
  TBUFX2 \read_data_2_tri[23]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[23]) );
  TBUFX2 \read_data_2_tri[22]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[22]) );
  TBUFX2 \read_data_2_tri[21]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[21]) );
  TBUFX2 \read_data_2_tri[20]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[20]) );
  TBUFX2 \read_data_2_tri[19]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[19]) );
  TBUFX2 \read_data_2_tri[18]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[18]) );
  TBUFX2 \read_data_2_tri[17]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[17]) );
  TBUFX2 \read_data_2_tri[16]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[16]) );
  TBUFX2 \read_data_2_tri[15]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[15]) );
  TBUFX2 \read_data_2_tri[14]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[14]) );
  TBUFX2 \read_data_2_tri[13]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[13]) );
  TBUFX2 \read_data_2_tri[12]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[12]) );
  TBUFX2 \read_data_2_tri[11]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[11]) );
  TBUFX2 \read_data_2_tri[10]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[10]) );
  TBUFX2 \read_data_2_tri[9]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[9]) );
  TBUFX2 \read_data_2_tri[8]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[8]) );
  TBUFX2 \read_data_2_tri[7]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[7]) );
  TBUFX2 \read_data_2_tri[6]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[6]) );
  TBUFX2 \read_data_2_tri[5]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[5]) );
  TBUFX2 \read_data_2_tri[3]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[3]) );
  TBUFX2 \read_data_2_tri[2]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[2]) );
  TBUFX2 \read_data_2_tri[1]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[1]) );
  TBUFX2 \read_data_2_tri[0]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[0]) );
  TBUFX2 \read_data_2_tri[4]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[4]) );
  TBUFX2 \read_data_2_tri[29]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[29]) );
  TBUFX2 \read_data_1_tri[9]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[9]) );
endmodule


module Register_File_WIDTH32_DEPTH5_0 ( clk, reset, read_enable_1, 
        read_enable_2, write_enable, read_index_1, read_index_2, write_index, 
        write_data, read_data_1, read_data_2 );
  input [4:0] read_index_1;
  input [4:0] read_index_2;
  input [4:0] write_index;
  input [31:0] write_data;
  output [31:0] read_data_1;
  output [31:0] read_data_2;
  input clk, reset, read_enable_1, read_enable_2, write_enable;

  tri   [31:0] read_data_1;
  tri   [31:0] read_data_2;

  TBUFX2 \read_data_1_tri[31]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[31]) );
  TBUFX2 \read_data_1_tri[30]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[30]) );
  TBUFX2 \read_data_1_tri[29]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[29]) );
  TBUFX2 \read_data_1_tri[28]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[28]) );
  TBUFX2 \read_data_1_tri[27]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[27]) );
  TBUFX2 \read_data_1_tri[26]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[26]) );
  TBUFX2 \read_data_1_tri[25]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[25]) );
  TBUFX2 \read_data_1_tri[24]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[24]) );
  TBUFX2 \read_data_1_tri[23]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[23]) );
  TBUFX2 \read_data_1_tri[22]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[22]) );
  TBUFX2 \read_data_1_tri[21]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[21]) );
  TBUFX2 \read_data_1_tri[20]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[20]) );
  TBUFX2 \read_data_1_tri[19]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[19]) );
  TBUFX2 \read_data_1_tri[18]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[18]) );
  TBUFX2 \read_data_1_tri[17]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[17]) );
  TBUFX2 \read_data_1_tri[16]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[16]) );
  TBUFX2 \read_data_1_tri[15]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[15]) );
  TBUFX2 \read_data_1_tri[14]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[14]) );
  TBUFX2 \read_data_1_tri[13]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[13]) );
  TBUFX2 \read_data_1_tri[12]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[12]) );
  TBUFX2 \read_data_1_tri[11]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[11]) );
  TBUFX2 \read_data_1_tri[10]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[10]) );
  TBUFX2 \read_data_1_tri[9]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[9]) );
  TBUFX2 \read_data_1_tri[8]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[8]) );
  TBUFX2 \read_data_1_tri[7]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[7]) );
  TBUFX2 \read_data_1_tri[6]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[6]) );
  TBUFX2 \read_data_1_tri[5]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[5]) );
  TBUFX2 \read_data_1_tri[4]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[4]) );
  TBUFX2 \read_data_1_tri[3]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[3]) );
  TBUFX2 \read_data_1_tri[2]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[2]) );
  TBUFX2 \read_data_1_tri[1]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[1]) );
  TBUFX2 \read_data_1_tri[0]  ( .A(1'b1), .EN(1'b0), .Y(read_data_1[0]) );
  TBUFX2 \read_data_2_tri[31]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[31]) );
  TBUFX2 \read_data_2_tri[30]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[30]) );
  TBUFX2 \read_data_2_tri[29]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[29]) );
  TBUFX2 \read_data_2_tri[28]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[28]) );
  TBUFX2 \read_data_2_tri[27]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[27]) );
  TBUFX2 \read_data_2_tri[26]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[26]) );
  TBUFX2 \read_data_2_tri[25]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[25]) );
  TBUFX2 \read_data_2_tri[24]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[24]) );
  TBUFX2 \read_data_2_tri[23]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[23]) );
  TBUFX2 \read_data_2_tri[22]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[22]) );
  TBUFX2 \read_data_2_tri[21]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[21]) );
  TBUFX2 \read_data_2_tri[20]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[20]) );
  TBUFX2 \read_data_2_tri[19]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[19]) );
  TBUFX2 \read_data_2_tri[18]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[18]) );
  TBUFX2 \read_data_2_tri[17]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[17]) );
  TBUFX2 \read_data_2_tri[16]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[16]) );
  TBUFX2 \read_data_2_tri[15]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[15]) );
  TBUFX2 \read_data_2_tri[14]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[14]) );
  TBUFX2 \read_data_2_tri[13]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[13]) );
  TBUFX2 \read_data_2_tri[12]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[12]) );
  TBUFX2 \read_data_2_tri[11]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[11]) );
  TBUFX2 \read_data_2_tri[10]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[10]) );
  TBUFX2 \read_data_2_tri[9]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[9]) );
  TBUFX2 \read_data_2_tri[8]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[8]) );
  TBUFX2 \read_data_2_tri[7]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[7]) );
  TBUFX2 \read_data_2_tri[6]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[6]) );
  TBUFX2 \read_data_2_tri[5]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[5]) );
  TBUFX2 \read_data_2_tri[4]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[4]) );
  TBUFX2 \read_data_2_tri[3]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[3]) );
  TBUFX2 \read_data_2_tri[2]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[2]) );
  TBUFX2 \read_data_2_tri[1]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[1]) );
  TBUFX2 \read_data_2_tri[0]  ( .A(1'b1), .EN(1'b0), .Y(read_data_2[0]) );
endmodule


module LUMOS ( clk, reset, trap, memoryData, memoryReady, memoryEnable, 
        memoryReadWrite, memoryAddress );
  inout [31:0] memoryData;
  output [31:0] memoryAddress;
  input clk, reset, memoryReady;
  output trap, memoryEnable, memoryReadWrite;
  wire   aluZeroRegister, aluSignRegister, N466, N467, N719, N721, N924, N965,
         N966, N968, N969, N971, N972, N1116, N1117, N1119, N1120, N1122,
         N1123, N1125, N1126, N1128, N1129, N1131, N1132, N1134, N1135, N1137,
         N1138, N1140, N1141, N1143, N1144, N1146, N1147, N1149, N1150, N1152,
         N1153, N1155, N1156, N1158, N1159, N1161, N1162, N1164, N1165, N1167,
         N1168, N1170, N1171, N1173, N1174, N1176, N1177, N1179, N1180, N1182,
         N1183, N1185, N1186, N1188, N1189, N1191, N1192, N1194, N1195, N1197,
         N1198, N1200, N1201, N1203, N1204, N1206, N1207, N1209, N1210,
         \arithmetic_logic_unit/N300 , \arithmetic_logic_unit/N298 ,
         \arithmetic_logic_unit/N294 , \arithmetic_logic_unit/N289 ,
         \arithmetic_logic_unit/N288 , \arithmetic_logic_unit/N286 ,
         \arithmetic_logic_unit/N284 , \arithmetic_logic_unit/N279 ,
         \arithmetic_logic_unit/N278 , \arithmetic_logic_unit/N277 ,
         \arithmetic_logic_unit/N276 , \arithmetic_logic_unit/N275 ,
         \arithmetic_logic_unit/N274 , \arithmetic_logic_unit/N273 ,
         \arithmetic_logic_unit/N272 , \arithmetic_logic_unit/N268 ,
         \arithmetic_logic_unit/N266 , \arithmetic_logic_unit/N151 ,
         \arithmetic_logic_unit/N150 , \arithmetic_logic_unit/N149 ,
         \arithmetic_logic_unit/N148 , \arithmetic_logic_unit/N147 ,
         \arithmetic_logic_unit/N146 , \arithmetic_logic_unit/N145 ,
         \arithmetic_logic_unit/N144 , \arithmetic_logic_unit/N143 ,
         \arithmetic_logic_unit/N142 , \arithmetic_logic_unit/N138 ,
         \arithmetic_logic_unit/N136 , \arithmetic_logic_unit/N132 ,
         \arithmetic_logic_unit/N127 , \arithmetic_logic_unit/N126 ,
         \arithmetic_logic_unit/N124 , \arithmetic_logic_unit/N122 ,
         \arithmetic_logic_unit/N119 , \arithmetic_logic_unit/N118 ,
         \arithmetic_logic_unit/N117 , \arithmetic_logic_unit/N116 ,
         \arithmetic_logic_unit/N115 , \arithmetic_logic_unit/N114 ,
         \arithmetic_logic_unit/N113 , \arithmetic_logic_unit/N112 ,
         \arithmetic_logic_unit/N111 , \arithmetic_logic_unit/N110 ,
         \arithmetic_logic_unit/N106 , \arithmetic_logic_unit/N104 ,
         \arithmetic_logic_unit/N100 , \arithmetic_logic_unit/N95 ,
         \arithmetic_logic_unit/N94 , \arithmetic_logic_unit/N92 ,
         \arithmetic_logic_unit/N90 , n61, n138, n217, n245, n504, n513, n515,
         n517, n518, n524, n526, n533, n535, n537, n538, n539, n540, n541,
         n542, n543, n544, n547, n549, n551, n553, n555, n557, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n627,
         n629, n631, n633, n635, n637, n639, n641, n643, n645, n647, n649,
         n651, n653, n655, n657, n659, n661, n663, n665, n667, n669, n671,
         n673, n675, n677, n679, n681, n683, n685, n847, n848, n849, n851,
         n853, n855, n871, n873, n875, n877, n879, n881, n883, n885, n887,
         n889, n891, n893, n895, n897, n899, n901, n903, n905, n907, n913,
         n917, n921, n923, n925, n927, n929, n931, n933, n941, n945, n947,
         n953, n955, n957, n959, n961, n963, n965, n967, n971, n977, n978,
         n980, n981, n982, n987, n989, n991, n993, n995, n996, n998, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1156, n1157, n1158, n1159, n1160, n1188, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1247, n1275, n1277, n1279, n1281, n1283, n1286, n1287, n1288, n1289,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1381, n1424, n1426, n1427, n1430, n1449, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1554,
         \ashr_1100_6/SH[3] , \ashr_1100_6/SH[2] , \ashr_1100_6/SH[1] ,
         \ashr_1100_6/SH[0] , \lt_x_1100_4/B[31] , \lt_x_1100_4/B[30] ,
         \lt_x_1100_4/B[29] , \lt_x_1100_4/B[28] , \lt_x_1100_4/B[27] ,
         \lt_x_1100_4/B[26] , \lt_x_1100_4/B[25] , \lt_x_1100_4/B[24] ,
         \lt_x_1100_4/B[23] , \lt_x_1100_4/B[22] , \lt_x_1100_4/B[21] ,
         \lt_x_1100_4/B[20] , \lt_x_1100_4/B[19] , \lt_x_1100_4/B[18] ,
         \lt_x_1100_4/B[17] , \lt_x_1100_4/B[16] , \lt_x_1100_4/B[15] ,
         \lt_x_1100_4/B[13] , \lt_x_1100_4/B[12] , \lt_x_1100_4/B[11] ,
         \lt_x_1100_4/B[10] , \lt_x_1100_4/B[9] , \lt_x_1100_4/B[8] ,
         \lt_x_1100_4/B[7] , \lt_x_1100_4/B[6] , \lt_x_1100_4/B[5] ,
         \sub_x_1100_2/A[31] , \sub_x_1100_2/A[30] , \sub_x_1100_2/A[29] ,
         \sub_x_1100_2/A[28] , \sub_x_1100_2/A[27] , \sub_x_1100_2/A[14] ,
         \sub_x_1100_2/A[13] , \sub_x_1100_2/A[12] , \sub_x_1100_2/A[11] ,
         \sub_x_1100_2/A[10] , \sub_x_1100_2/A[8] , \sub_x_1100_2/A[7] ,
         \sub_x_1100_2/A[6] , \sub_x_1100_2/A[5] , \sub_x_1100_2/A[4] ,
         \sub_x_1100_2/A[2] , \sub_x_1100_2/A[0] , \sub_x_1100_2/B[4] ,
         \sub_x_1100_2/n228 , \sub_x_1100_2/n227 , \sub_x_1100_2/n216 ,
         \sub_x_1100_2/n198 , \sub_x_1100_2/n174 , \sub_x_1100_2/n170 ,
         \sub_x_1100_2/n169 , \sub_x_1100_2/n166 , \sub_x_1100_2/n163 ,
         \sub_x_1100_2/n161 , \sub_x_1100_2/n160 , \sub_x_1100_2/n155 ,
         \sub_x_1100_2/n152 , \sub_x_1100_2/n150 , \sub_x_1100_2/n144 ,
         \sub_x_1100_2/n142 , \sub_x_1100_2/n139 , \sub_x_1100_2/n133 ,
         \sub_x_1100_2/n131 , \sub_x_1100_2/n129 , \sub_x_1100_2/n124 ,
         \sub_x_1100_2/n121 , \sub_x_1100_2/n119 , \sub_x_1100_2/n117 ,
         \sub_x_1100_2/n116 , \sub_x_1100_2/n108 , \sub_x_1100_2/n106 ,
         \sub_x_1100_2/n104 , \sub_x_1100_2/n99 , \sub_x_1100_2/n96 ,
         \sub_x_1100_2/n94 , \sub_x_1100_2/n92 , \sub_x_1100_2/n90 ,
         \sub_x_1100_2/n89 , \sub_x_1100_2/n84 , \sub_x_1100_2/n79 ,
         \sub_x_1100_2/n77 , \sub_x_1100_2/n72 , \sub_x_1100_2/n69 ,
         \sub_x_1100_2/n64 , \sub_x_1100_2/n53 , \sub_x_1100_2/n37 ,
         \sub_x_1100_2/n31 , \sub_x_1100_2/n30 , \add_x_1100_1/n197 ,
         \add_x_1100_1/n195 , \add_x_1100_1/n193 , \add_x_1100_1/n192 ,
         \add_x_1100_1/n188 , \add_x_1100_1/n187 , \add_x_1100_1/n186 ,
         \add_x_1100_1/n166 , \add_x_1100_1/n165 , \add_x_1100_1/n162 ,
         \add_x_1100_1/n159 , \add_x_1100_1/n157 , \add_x_1100_1/n156 ,
         \add_x_1100_1/n151 , \add_x_1100_1/n148 , \add_x_1100_1/n146 ,
         \add_x_1100_1/n140 , \add_x_1100_1/n138 , \add_x_1100_1/n136 ,
         \add_x_1100_1/n135 , \add_x_1100_1/n129 , \add_x_1100_1/n127 ,
         \add_x_1100_1/n126 , \add_x_1100_1/n125 , \add_x_1100_1/n120 ,
         \add_x_1100_1/n117 , \add_x_1100_1/n115 , \add_x_1100_1/n113 ,
         \add_x_1100_1/n112 , \add_x_1100_1/n104 , \add_x_1100_1/n102 ,
         \add_x_1100_1/n100 , \add_x_1100_1/n96 , \add_x_1100_1/n95 ,
         \add_x_1100_1/n92 , \add_x_1100_1/n90 , \add_x_1100_1/n88 ,
         \add_x_1100_1/n86 , \add_x_1100_1/n85 , \add_x_1100_1/n80 ,
         \add_x_1100_1/n75 , \add_x_1100_1/n73 , \add_x_1100_1/n68 ,
         \add_x_1100_1/n65 , \add_x_1100_1/n49 , \add_x_1100_1/n33 ,
         \add_x_1100_1/n32 , \add_x_1100_1/n31 , \add_x_1100_1/n30 ,
         \sub_x_1100_2/n32 , n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375;
  wire   [31:0] pc;
  wire   [31:0] memoryDataRegister;
  wire   [31:0] RS2;
  wire   [31:0] RS1;
  wire   [31:0] aluOperand1;
  wire   [31:0] aluResultRegister;
  tri   clk;
  tri   reset;
  tri   [31:0] memoryData;
  tri   memoryReadWrite;
  tri   [24:15] ir;
  tri   ir_11;
  tri   ir_10;
  tri   ir_9;
  tri   ir_8;
  tri   ir_7;
  tri   [6:0] opcode;
  tri   [2:0] funct3;
  tri   [6:0] funct7;
  tri   [4:0] nextState;
  tri   fpuReady;
  tri   pcWrite;
  tri   irWrite;
  tri   [3:0] aluOperation;
  tri   [1:0] aluSrcA;
  tri   [1:0] aluSrcB;
  tri   instructionOrData;
  tri   [2:0] instructionType;
  tri   [1:0] fpuOperation;
  tri   [31:0] aluResult;
  tri   [31:0] FRS2;
  tri   [31:0] readData1;
  tri   [31:0] readData2;
  tri   [31:0] fpuResult;
  tri   [31:0] fixedPointReadData1;
  tri   [31:0] fixedPointReadData2;
  tri   [31:0] FRS1;
  tri   [31:0] immediate;
  tri   \opcode[1] ;
  tri   \opcode[0] ;
  tri   \funct3[0] ;
  assign trap = 1'b1;

  Register_File_WIDTH32_DEPTH5_1 register_file ( .clk(1'b0), .reset(1'b0), 
        .read_enable_1(1'b1), .read_enable_2(1'b1), .write_enable(1'b0), 
        .read_index_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .read_index_2({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .write_index({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .write_data({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .read_data_1(readData1), .read_data_2(readData2) );
  Register_File_WIDTH32_DEPTH5_0 fixed_point_register_file ( .clk(1'b0), 
        .reset(1'b0), .read_enable_1(1'b1), .read_enable_2(1'b1), 
        .write_enable(1'b0), .read_index_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .read_index_2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .write_index({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .write_data({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .read_data_1(fixedPointReadData1), .read_data_2(
        fixedPointReadData2) );
  Fixed_Point_Unit fixed_point_unit ( .clk(clk), .reset(reset), .operand_1(
        FRS1), .operand_2(FRS2), .operation(fpuOperation), .result(fpuResult), 
        .ready(fpuReady) );
  DFFPOSX1 aluSignRegister_reg ( .D(n1850), .CLK(clk), .Q(aluSignRegister) );
  DFFPOSX1 \pc_reg[0]  ( .D(n1458), .CLK(clk), .Q(pc[0]) );
  DFFPOSX1 \RS1_reg[31]  ( .D(readData1[31]), .CLK(clk), .Q(RS1[31]) );
  DFFPOSX1 aluZeroRegister_reg ( .D(n1554), .CLK(clk), .Q(aluZeroRegister) );
  DFFSR \state_reg[1]  ( .D(n998), .CLK(clk), .R(1'b1), .S(n4364), .Q(n1000)
         );
  DFFSR \state_reg[2]  ( .D(n996), .CLK(clk), .R(1'b1), .S(n4364), .Q(n1104)
         );
  DFFSR \state_reg[3]  ( .D(n993), .CLK(clk), .R(1'b1), .S(n4364), .Q(n995) );
  DFFPOSX1 \FRS1_reg[31]  ( .D(fixedPointReadData1[31]), .CLK(clk), .Q(
        FRS1[31]) );
  DFFPOSX1 \RS1_reg[30]  ( .D(readData1[30]), .CLK(clk), .Q(RS1[30]) );
  DFFPOSX1 \RS1_reg[29]  ( .D(readData1[29]), .CLK(clk), .Q(RS1[29]) );
  DFFPOSX1 \RS1_reg[28]  ( .D(readData1[28]), .CLK(clk), .Q(RS1[28]) );
  DFFPOSX1 \RS1_reg[27]  ( .D(readData1[27]), .CLK(clk), .Q(RS1[27]) );
  DFFPOSX1 \RS1_reg[26]  ( .D(readData1[26]), .CLK(clk), .Q(RS1[26]) );
  DFFPOSX1 \RS1_reg[25]  ( .D(readData1[25]), .CLK(clk), .Q(RS1[25]) );
  DFFPOSX1 \RS1_reg[24]  ( .D(readData1[24]), .CLK(clk), .Q(RS1[24]) );
  DFFPOSX1 \RS1_reg[23]  ( .D(readData1[23]), .CLK(clk), .Q(RS1[23]) );
  DFFPOSX1 \RS1_reg[22]  ( .D(readData1[22]), .CLK(clk), .Q(RS1[22]) );
  DFFPOSX1 \RS1_reg[21]  ( .D(readData1[21]), .CLK(clk), .Q(RS1[21]) );
  DFFPOSX1 \RS1_reg[20]  ( .D(readData1[20]), .CLK(clk), .Q(RS1[20]) );
  DFFPOSX1 \RS1_reg[19]  ( .D(readData1[19]), .CLK(clk), .Q(RS1[19]) );
  DFFPOSX1 \RS1_reg[18]  ( .D(readData1[18]), .CLK(clk), .Q(RS1[18]) );
  DFFPOSX1 \RS1_reg[17]  ( .D(readData1[17]), .CLK(clk), .Q(RS1[17]) );
  DFFPOSX1 \RS1_reg[16]  ( .D(readData1[16]), .CLK(clk), .Q(RS1[16]) );
  DFFPOSX1 \RS1_reg[15]  ( .D(readData1[15]), .CLK(clk), .Q(RS1[15]) );
  DFFPOSX1 \RS1_reg[14]  ( .D(readData1[14]), .CLK(clk), .Q(RS1[14]) );
  DFFPOSX1 \RS1_reg[13]  ( .D(readData1[13]), .CLK(clk), .Q(RS1[13]) );
  DFFPOSX1 \RS1_reg[12]  ( .D(readData1[12]), .CLK(clk), .Q(RS1[12]) );
  DFFPOSX1 \RS1_reg[11]  ( .D(readData1[11]), .CLK(clk), .Q(RS1[11]) );
  DFFPOSX1 \RS1_reg[10]  ( .D(readData1[10]), .CLK(clk), .Q(RS1[10]) );
  DFFPOSX1 \RS1_reg[9]  ( .D(readData1[9]), .CLK(clk), .Q(RS1[9]) );
  DFFPOSX1 \RS1_reg[8]  ( .D(readData1[8]), .CLK(clk), .Q(RS1[8]) );
  DFFPOSX1 \RS1_reg[7]  ( .D(readData1[7]), .CLK(clk), .Q(RS1[7]) );
  DFFPOSX1 \RS1_reg[6]  ( .D(readData1[6]), .CLK(clk), .Q(RS1[6]) );
  DFFPOSX1 \RS1_reg[5]  ( .D(readData1[5]), .CLK(clk), .Q(RS1[5]) );
  DFFPOSX1 \RS1_reg[4]  ( .D(readData1[4]), .CLK(clk), .Q(RS1[4]) );
  DFFPOSX1 \RS1_reg[3]  ( .D(readData1[3]), .CLK(clk), .Q(RS1[3]) );
  DFFPOSX1 \RS1_reg[2]  ( .D(readData1[2]), .CLK(clk), .Q(RS1[2]) );
  DFFPOSX1 \RS1_reg[1]  ( .D(readData1[1]), .CLK(clk), .Q(RS1[1]) );
  DFFPOSX1 \RS1_reg[0]  ( .D(readData1[0]), .CLK(clk), .Q(RS1[0]) );
  DFFPOSX1 \RS2_reg[31]  ( .D(readData2[31]), .CLK(clk), .Q(RS2[31]) );
  DFFPOSX1 \RS2_reg[30]  ( .D(readData2[30]), .CLK(clk), .Q(RS2[30]) );
  DFFPOSX1 \RS2_reg[29]  ( .D(readData2[29]), .CLK(clk), .Q(RS2[29]) );
  DFFPOSX1 \RS2_reg[28]  ( .D(readData2[28]), .CLK(clk), .Q(RS2[28]) );
  DFFPOSX1 \RS2_reg[27]  ( .D(readData2[27]), .CLK(clk), .Q(RS2[27]) );
  DFFPOSX1 \RS2_reg[26]  ( .D(readData2[26]), .CLK(clk), .Q(RS2[26]) );
  DFFPOSX1 \RS2_reg[25]  ( .D(readData2[25]), .CLK(clk), .Q(RS2[25]) );
  DFFPOSX1 \RS2_reg[24]  ( .D(readData2[24]), .CLK(clk), .Q(RS2[24]) );
  DFFPOSX1 \RS2_reg[23]  ( .D(readData2[23]), .CLK(clk), .Q(RS2[23]) );
  DFFPOSX1 \RS2_reg[22]  ( .D(readData2[22]), .CLK(clk), .Q(RS2[22]) );
  DFFPOSX1 \RS2_reg[21]  ( .D(readData2[21]), .CLK(clk), .Q(RS2[21]) );
  DFFPOSX1 \RS2_reg[20]  ( .D(readData2[20]), .CLK(clk), .Q(RS2[20]) );
  DFFPOSX1 \RS2_reg[19]  ( .D(readData2[19]), .CLK(clk), .Q(RS2[19]) );
  DFFPOSX1 \RS2_reg[18]  ( .D(readData2[18]), .CLK(clk), .Q(RS2[18]) );
  DFFPOSX1 \RS2_reg[17]  ( .D(readData2[17]), .CLK(clk), .Q(RS2[17]) );
  DFFPOSX1 \RS2_reg[16]  ( .D(readData2[16]), .CLK(clk), .Q(RS2[16]) );
  DFFPOSX1 \RS2_reg[15]  ( .D(readData2[15]), .CLK(clk), .Q(RS2[15]) );
  DFFPOSX1 \RS2_reg[14]  ( .D(readData2[14]), .CLK(clk), .Q(RS2[14]) );
  DFFPOSX1 \RS2_reg[13]  ( .D(readData2[13]), .CLK(clk), .Q(RS2[13]) );
  DFFPOSX1 \RS2_reg[12]  ( .D(readData2[12]), .CLK(clk), .Q(RS2[12]) );
  DFFPOSX1 \RS2_reg[11]  ( .D(readData2[11]), .CLK(clk), .Q(RS2[11]) );
  DFFPOSX1 \RS2_reg[10]  ( .D(readData2[10]), .CLK(clk), .Q(RS2[10]) );
  DFFPOSX1 \RS2_reg[9]  ( .D(readData2[9]), .CLK(clk), .Q(RS2[9]) );
  DFFPOSX1 \RS2_reg[8]  ( .D(readData2[8]), .CLK(clk), .Q(RS2[8]) );
  DFFPOSX1 \RS2_reg[7]  ( .D(readData2[7]), .CLK(clk), .Q(RS2[7]) );
  DFFPOSX1 \RS2_reg[6]  ( .D(readData2[6]), .CLK(clk), .Q(RS2[6]) );
  DFFPOSX1 \RS2_reg[5]  ( .D(readData2[5]), .CLK(clk), .Q(RS2[5]) );
  DFFPOSX1 \RS2_reg[4]  ( .D(readData2[4]), .CLK(clk), .Q(RS2[4]) );
  DFFPOSX1 \RS2_reg[3]  ( .D(readData2[3]), .CLK(clk), .Q(RS2[3]) );
  DFFPOSX1 \RS2_reg[2]  ( .D(readData2[2]), .CLK(clk), .Q(RS2[2]) );
  DFFPOSX1 \RS2_reg[1]  ( .D(readData2[1]), .CLK(clk), .Q(RS2[1]) );
  DFFPOSX1 \RS2_reg[0]  ( .D(readData2[0]), .CLK(clk), .Q(RS2[0]) );
  DFFPOSX1 \FRS1_reg[30]  ( .D(fixedPointReadData1[30]), .CLK(clk), .Q(
        FRS1[30]) );
  DFFPOSX1 \FRS1_reg[29]  ( .D(fixedPointReadData1[29]), .CLK(clk), .Q(
        FRS1[29]) );
  DFFPOSX1 \FRS1_reg[28]  ( .D(fixedPointReadData1[28]), .CLK(clk), .Q(
        FRS1[28]) );
  DFFPOSX1 \FRS1_reg[27]  ( .D(fixedPointReadData1[27]), .CLK(clk), .Q(
        FRS1[27]) );
  DFFPOSX1 \FRS1_reg[26]  ( .D(fixedPointReadData1[26]), .CLK(clk), .Q(
        FRS1[26]) );
  DFFPOSX1 \FRS1_reg[25]  ( .D(fixedPointReadData1[25]), .CLK(clk), .Q(
        FRS1[25]) );
  DFFPOSX1 \FRS1_reg[24]  ( .D(fixedPointReadData1[24]), .CLK(clk), .Q(
        FRS1[24]) );
  DFFPOSX1 \FRS1_reg[23]  ( .D(fixedPointReadData1[23]), .CLK(clk), .Q(
        FRS1[23]) );
  DFFPOSX1 \FRS1_reg[22]  ( .D(fixedPointReadData1[22]), .CLK(clk), .Q(
        FRS1[22]) );
  DFFPOSX1 \FRS1_reg[21]  ( .D(fixedPointReadData1[21]), .CLK(clk), .Q(
        FRS1[21]) );
  DFFPOSX1 \FRS1_reg[20]  ( .D(fixedPointReadData1[20]), .CLK(clk), .Q(
        FRS1[20]) );
  DFFPOSX1 \FRS1_reg[19]  ( .D(fixedPointReadData1[19]), .CLK(clk), .Q(
        FRS1[19]) );
  DFFPOSX1 \FRS1_reg[18]  ( .D(fixedPointReadData1[18]), .CLK(clk), .Q(
        FRS1[18]) );
  DFFPOSX1 \FRS1_reg[17]  ( .D(fixedPointReadData1[17]), .CLK(clk), .Q(
        FRS1[17]) );
  DFFPOSX1 \FRS1_reg[16]  ( .D(fixedPointReadData1[16]), .CLK(clk), .Q(
        FRS1[16]) );
  DFFPOSX1 \FRS1_reg[15]  ( .D(fixedPointReadData1[15]), .CLK(clk), .Q(
        FRS1[15]) );
  DFFPOSX1 \FRS1_reg[14]  ( .D(fixedPointReadData1[14]), .CLK(clk), .Q(
        FRS1[14]) );
  DFFPOSX1 \FRS1_reg[13]  ( .D(fixedPointReadData1[13]), .CLK(clk), .Q(
        FRS1[13]) );
  DFFPOSX1 \FRS1_reg[12]  ( .D(fixedPointReadData1[12]), .CLK(clk), .Q(
        FRS1[12]) );
  DFFPOSX1 \FRS1_reg[11]  ( .D(fixedPointReadData1[11]), .CLK(clk), .Q(
        FRS1[11]) );
  DFFPOSX1 \FRS1_reg[10]  ( .D(fixedPointReadData1[10]), .CLK(clk), .Q(
        FRS1[10]) );
  DFFPOSX1 \FRS1_reg[9]  ( .D(fixedPointReadData1[9]), .CLK(clk), .Q(FRS1[9])
         );
  DFFPOSX1 \FRS1_reg[8]  ( .D(fixedPointReadData1[8]), .CLK(clk), .Q(FRS1[8])
         );
  DFFPOSX1 \FRS1_reg[7]  ( .D(fixedPointReadData1[7]), .CLK(clk), .Q(FRS1[7])
         );
  DFFPOSX1 \FRS1_reg[6]  ( .D(fixedPointReadData1[6]), .CLK(clk), .Q(FRS1[6])
         );
  DFFPOSX1 \FRS1_reg[5]  ( .D(fixedPointReadData1[5]), .CLK(clk), .Q(FRS1[5])
         );
  DFFPOSX1 \FRS1_reg[4]  ( .D(fixedPointReadData1[4]), .CLK(clk), .Q(FRS1[4])
         );
  DFFPOSX1 \FRS1_reg[3]  ( .D(fixedPointReadData1[3]), .CLK(clk), .Q(FRS1[3])
         );
  DFFPOSX1 \FRS1_reg[2]  ( .D(fixedPointReadData1[2]), .CLK(clk), .Q(FRS1[2])
         );
  DFFPOSX1 \FRS1_reg[1]  ( .D(fixedPointReadData1[1]), .CLK(clk), .Q(FRS1[1])
         );
  DFFPOSX1 \FRS1_reg[0]  ( .D(fixedPointReadData1[0]), .CLK(clk), .Q(FRS1[0])
         );
  DFFPOSX1 \FRS2_reg[31]  ( .D(fixedPointReadData2[31]), .CLK(clk), .Q(
        FRS2[31]) );
  DFFPOSX1 \FRS2_reg[30]  ( .D(fixedPointReadData2[30]), .CLK(clk), .Q(
        FRS2[30]) );
  DFFPOSX1 \FRS2_reg[29]  ( .D(fixedPointReadData2[29]), .CLK(clk), .Q(
        FRS2[29]) );
  DFFPOSX1 \FRS2_reg[28]  ( .D(fixedPointReadData2[28]), .CLK(clk), .Q(
        FRS2[28]) );
  DFFPOSX1 \FRS2_reg[27]  ( .D(fixedPointReadData2[27]), .CLK(clk), .Q(
        FRS2[27]) );
  DFFPOSX1 \FRS2_reg[26]  ( .D(fixedPointReadData2[26]), .CLK(clk), .Q(
        FRS2[26]) );
  DFFPOSX1 \FRS2_reg[25]  ( .D(fixedPointReadData2[25]), .CLK(clk), .Q(
        FRS2[25]) );
  DFFPOSX1 \FRS2_reg[24]  ( .D(fixedPointReadData2[24]), .CLK(clk), .Q(
        FRS2[24]) );
  DFFPOSX1 \FRS2_reg[23]  ( .D(fixedPointReadData2[23]), .CLK(clk), .Q(
        FRS2[23]) );
  DFFPOSX1 \FRS2_reg[22]  ( .D(fixedPointReadData2[22]), .CLK(clk), .Q(
        FRS2[22]) );
  DFFPOSX1 \FRS2_reg[21]  ( .D(fixedPointReadData2[21]), .CLK(clk), .Q(
        FRS2[21]) );
  DFFPOSX1 \FRS2_reg[20]  ( .D(fixedPointReadData2[20]), .CLK(clk), .Q(
        FRS2[20]) );
  DFFPOSX1 \FRS2_reg[19]  ( .D(fixedPointReadData2[19]), .CLK(clk), .Q(
        FRS2[19]) );
  DFFPOSX1 \FRS2_reg[18]  ( .D(fixedPointReadData2[18]), .CLK(clk), .Q(
        FRS2[18]) );
  DFFPOSX1 \FRS2_reg[17]  ( .D(fixedPointReadData2[17]), .CLK(clk), .Q(
        FRS2[17]) );
  DFFPOSX1 \FRS2_reg[16]  ( .D(fixedPointReadData2[16]), .CLK(clk), .Q(
        FRS2[16]) );
  DFFPOSX1 \FRS2_reg[15]  ( .D(fixedPointReadData2[15]), .CLK(clk), .Q(
        FRS2[15]) );
  DFFPOSX1 \FRS2_reg[14]  ( .D(fixedPointReadData2[14]), .CLK(clk), .Q(
        FRS2[14]) );
  DFFPOSX1 \FRS2_reg[13]  ( .D(fixedPointReadData2[13]), .CLK(clk), .Q(
        FRS2[13]) );
  DFFPOSX1 \FRS2_reg[12]  ( .D(fixedPointReadData2[12]), .CLK(clk), .Q(
        FRS2[12]) );
  DFFPOSX1 \FRS2_reg[11]  ( .D(fixedPointReadData2[11]), .CLK(clk), .Q(
        FRS2[11]) );
  DFFPOSX1 \FRS2_reg[10]  ( .D(fixedPointReadData2[10]), .CLK(clk), .Q(
        FRS2[10]) );
  DFFPOSX1 \FRS2_reg[9]  ( .D(fixedPointReadData2[9]), .CLK(clk), .Q(FRS2[9])
         );
  DFFPOSX1 \FRS2_reg[8]  ( .D(fixedPointReadData2[8]), .CLK(clk), .Q(FRS2[8])
         );
  DFFPOSX1 \FRS2_reg[7]  ( .D(fixedPointReadData2[7]), .CLK(clk), .Q(FRS2[7])
         );
  DFFPOSX1 \FRS2_reg[6]  ( .D(fixedPointReadData2[6]), .CLK(clk), .Q(FRS2[6])
         );
  DFFPOSX1 \FRS2_reg[5]  ( .D(fixedPointReadData2[5]), .CLK(clk), .Q(FRS2[5])
         );
  DFFPOSX1 \FRS2_reg[4]  ( .D(fixedPointReadData2[4]), .CLK(clk), .Q(FRS2[4])
         );
  DFFPOSX1 \FRS2_reg[3]  ( .D(fixedPointReadData2[3]), .CLK(clk), .Q(FRS2[3])
         );
  DFFPOSX1 \FRS2_reg[2]  ( .D(fixedPointReadData2[2]), .CLK(clk), .Q(FRS2[2])
         );
  DFFPOSX1 \FRS2_reg[1]  ( .D(fixedPointReadData2[1]), .CLK(clk), .Q(FRS2[1])
         );
  DFFPOSX1 \FRS2_reg[0]  ( .D(fixedPointReadData2[0]), .CLK(clk), .Q(FRS2[0])
         );
  DFFPOSX1 \memoryDataRegister_reg[0]  ( .D(n2506), .CLK(clk), .Q(
        memoryDataRegister[0]) );
  DFFPOSX1 \ir_reg[0]  ( .D(n1017), .CLK(clk), .Q(N1209) );
  DFFPOSX1 \memoryDataRegister_reg[2]  ( .D(n2510), .CLK(clk), .Q(
        memoryDataRegister[2]) );
  DFFPOSX1 \ir_reg[2]  ( .D(n1016), .CLK(clk), .Q(N1203) );
  DFFSR \state_reg[0]  ( .D(n991), .CLK(clk), .R(1'b1), .S(n4364), .Q(n987) );
  LATCH memoryEnable_reg ( .CLK(n3054), .D(n3154), .Q(memoryEnable) );
  DFFPOSX1 \ir_reg[14]  ( .D(n1010), .CLK(clk), .Q(N1167) );
  DFFSR \state_reg[4]  ( .D(n989), .CLK(clk), .R(1'b1), .S(n4364), .Q(n1103)
         );
  DFFPOSX1 \ir_tri_enable_reg[31]  ( .D(n2630), .CLK(clk), .Q(N1117) );
  DFFPOSX1 \ir_tri_enable_reg[30]  ( .D(n2628), .CLK(clk), .Q(N1120) );
  DFFPOSX1 \ir_tri_enable_reg[29]  ( .D(n2626), .CLK(clk), .Q(N1123) );
  DFFPOSX1 \ir_tri_enable_reg[28]  ( .D(n2624), .CLK(clk), .Q(N1126) );
  DFFPOSX1 \ir_tri_enable_reg[27]  ( .D(n2622), .CLK(clk), .Q(N1129) );
  DFFPOSX1 \ir_tri_enable_reg[26]  ( .D(n2620), .CLK(clk), .Q(N1132) );
  DFFPOSX1 \ir_tri_enable_reg[25]  ( .D(n2618), .CLK(clk), .Q(N1135) );
  DFFPOSX1 \ir_tri_enable_reg[24]  ( .D(n2616), .CLK(clk), .Q(N1138) );
  DFFPOSX1 \ir_tri_enable_reg[23]  ( .D(n2614), .CLK(clk), .Q(N1141) );
  DFFPOSX1 \ir_tri_enable_reg[22]  ( .D(n2612), .CLK(clk), .Q(N1144) );
  DFFPOSX1 \ir_tri_enable_reg[21]  ( .D(n2610), .CLK(clk), .Q(N1147) );
  DFFPOSX1 \ir_tri_enable_reg[20]  ( .D(n2608), .CLK(clk), .Q(N1150) );
  DFFPOSX1 \ir_tri_enable_reg[19]  ( .D(n2606), .CLK(clk), .Q(N1153) );
  DFFPOSX1 \ir_tri_enable_reg[18]  ( .D(n2604), .CLK(clk), .Q(N1156) );
  DFFPOSX1 \ir_tri_enable_reg[17]  ( .D(n2602), .CLK(clk), .Q(N1159) );
  DFFPOSX1 \ir_tri_enable_reg[16]  ( .D(n2600), .CLK(clk), .Q(N1162) );
  DFFPOSX1 \ir_tri_enable_reg[15]  ( .D(n2598), .CLK(clk), .Q(N1165) );
  DFFPOSX1 \ir_tri_enable_reg[14]  ( .D(n2596), .CLK(clk), .Q(N1168) );
  DFFPOSX1 \ir_tri_enable_reg[13]  ( .D(n2594), .CLK(clk), .Q(N1171) );
  DFFPOSX1 \ir_tri_enable_reg[12]  ( .D(n2592), .CLK(clk), .Q(N1174) );
  DFFPOSX1 \ir_tri_enable_reg[11]  ( .D(n2590), .CLK(clk), .Q(N1177) );
  DFFPOSX1 \ir_tri_enable_reg[10]  ( .D(n2588), .CLK(clk), .Q(N1180) );
  DFFPOSX1 \ir_tri_enable_reg[9]  ( .D(n2586), .CLK(clk), .Q(N1183) );
  DFFPOSX1 \ir_tri_enable_reg[8]  ( .D(n2584), .CLK(clk), .Q(N1186) );
  DFFPOSX1 \ir_tri_enable_reg[7]  ( .D(n2582), .CLK(clk), .Q(N1189) );
  DFFPOSX1 \ir_tri_enable_reg[6]  ( .D(n2580), .CLK(clk), .Q(N1192) );
  DFFPOSX1 \ir_tri_enable_reg[5]  ( .D(n2578), .CLK(clk), .Q(N1195) );
  DFFPOSX1 \ir_tri_enable_reg[4]  ( .D(n2576), .CLK(clk), .Q(N1198) );
  DFFPOSX1 \ir_tri_enable_reg[3]  ( .D(n2574), .CLK(clk), .Q(N1201) );
  DFFPOSX1 \ir_tri_enable_reg[2]  ( .D(n2572), .CLK(clk), .Q(N1204) );
  DFFPOSX1 \ir_tri_enable_reg[1]  ( .D(n2570), .CLK(clk), .Q(N1207) );
  DFFPOSX1 \ir_tri_enable_reg[0]  ( .D(n2568), .CLK(clk), .Q(N1210) );
  DFFPOSX1 \memoryDataRegister_reg[6]  ( .D(n2518), .CLK(clk), .Q(
        memoryDataRegister[6]) );
  DFFPOSX1 \ir_reg[6]  ( .D(n1014), .CLK(clk), .Q(N1191) );
  DFFPOSX1 \memoryDataRegister_reg[5]  ( .D(n2516), .CLK(clk), .Q(
        memoryDataRegister[5]) );
  DFFPOSX1 \ir_reg[5]  ( .D(n1020), .CLK(clk), .Q(N1194) );
  DFFPOSX1 \memoryDataRegister_reg[4]  ( .D(n2514), .CLK(clk), .Q(
        memoryDataRegister[4]) );
  DFFPOSX1 \ir_reg[4]  ( .D(n1015), .CLK(clk), .Q(N1197) );
  DFFPOSX1 \memoryDataRegister_reg[3]  ( .D(n2512), .CLK(clk), .Q(
        memoryDataRegister[3]) );
  DFFPOSX1 \ir_reg[3]  ( .D(n1019), .CLK(clk), .Q(N1200) );
  DFFPOSX1 \memoryDataRegister_reg[7]  ( .D(n2520), .CLK(clk), .Q(
        memoryDataRegister[7]) );
  DFFPOSX1 \ir_reg[7]  ( .D(n1021), .CLK(clk), .Q(N1188) );
  DFFPOSX1 \memoryDataRegister_reg[8]  ( .D(n2522), .CLK(clk), .Q(
        memoryDataRegister[8]) );
  DFFPOSX1 \ir_reg[8]  ( .D(n1013), .CLK(clk), .Q(N1185) );
  DFFPOSX1 \memoryDataRegister_reg[9]  ( .D(n2524), .CLK(clk), .Q(
        memoryDataRegister[9]) );
  DFFPOSX1 \ir_reg[9]  ( .D(n1022), .CLK(clk), .Q(N1182) );
  DFFPOSX1 \memoryDataRegister_reg[10]  ( .D(n2526), .CLK(clk), .Q(
        memoryDataRegister[10]) );
  DFFPOSX1 \ir_reg[10]  ( .D(n1012), .CLK(clk), .Q(N1179) );
  DFFPOSX1 \memoryDataRegister_reg[11]  ( .D(n2528), .CLK(clk), .Q(
        memoryDataRegister[11]) );
  DFFPOSX1 \ir_reg[11]  ( .D(n1023), .CLK(clk), .Q(N1176) );
  DFFPOSX1 \memoryDataRegister_reg[12]  ( .D(n2530), .CLK(clk), .Q(
        memoryDataRegister[12]) );
  DFFPOSX1 \ir_reg[12]  ( .D(n1011), .CLK(clk), .Q(N1173) );
  DFFPOSX1 \memoryDataRegister_reg[13]  ( .D(n2532), .CLK(clk), .Q(
        memoryDataRegister[13]) );
  DFFPOSX1 \ir_reg[13]  ( .D(n1024), .CLK(clk), .Q(N1170) );
  DFFPOSX1 \memoryDataRegister_reg[14]  ( .D(n2534), .CLK(clk), .Q(
        memoryDataRegister[14]) );
  DFFPOSX1 \memoryDataRegister_reg[15]  ( .D(n2536), .CLK(clk), .Q(
        memoryDataRegister[15]) );
  DFFPOSX1 \ir_reg[15]  ( .D(n1025), .CLK(clk), .Q(N1164) );
  DFFPOSX1 \memoryDataRegister_reg[17]  ( .D(n2540), .CLK(clk), .Q(
        memoryDataRegister[17]) );
  DFFPOSX1 \ir_reg[17]  ( .D(n1026), .CLK(clk), .Q(N1158) );
  DFFPOSX1 \memoryDataRegister_reg[19]  ( .D(n2544), .CLK(clk), .Q(
        memoryDataRegister[19]) );
  DFFPOSX1 \ir_reg[19]  ( .D(n1027), .CLK(clk), .Q(N1152) );
  DFFPOSX1 \memoryDataRegister_reg[21]  ( .D(n2548), .CLK(clk), .Q(
        memoryDataRegister[21]) );
  DFFPOSX1 \ir_reg[21]  ( .D(n1028), .CLK(clk), .Q(N1146) );
  DFFPOSX1 \memoryDataRegister_reg[23]  ( .D(n2552), .CLK(clk), .Q(
        memoryDataRegister[23]) );
  DFFPOSX1 \ir_reg[23]  ( .D(n1029), .CLK(clk), .Q(N1140) );
  DFFPOSX1 \memoryDataRegister_reg[25]  ( .D(n2556), .CLK(clk), .Q(
        memoryDataRegister[25]) );
  DFFPOSX1 \ir_reg[25]  ( .D(n1030), .CLK(clk), .Q(N1134) );
  DFFPOSX1 \memoryDataRegister_reg[27]  ( .D(n2560), .CLK(clk), .Q(
        memoryDataRegister[27]) );
  DFFPOSX1 \ir_reg[27]  ( .D(n1031), .CLK(clk), .Q(N1128) );
  DFFPOSX1 \memoryDataRegister_reg[29]  ( .D(n2564), .CLK(clk), .Q(
        memoryDataRegister[29]) );
  DFFPOSX1 \ir_reg[29]  ( .D(n1032), .CLK(clk), .Q(N1122) );
  LATCH \instructionType_reg[2]  ( .CLK(n4358), .D(N467), .Q(N965) );
  LATCH \instructionType_reg[0]  ( .CLK(n4358), .D(n2465), .Q(N971) );
  LATCH \instructionType_reg[1]  ( .CLK(n4358), .D(N466), .Q(N968) );
  DFFPOSX1 \memoryDataRegister_reg[16]  ( .D(n2538), .CLK(clk), .Q(
        memoryDataRegister[16]) );
  DFFPOSX1 \ir_reg[16]  ( .D(n1009), .CLK(clk), .Q(N1161) );
  DFFPOSX1 \memoryDataRegister_reg[18]  ( .D(n2542), .CLK(clk), .Q(
        memoryDataRegister[18]) );
  DFFPOSX1 \ir_reg[18]  ( .D(n1008), .CLK(clk), .Q(N1155) );
  DFFPOSX1 \memoryDataRegister_reg[20]  ( .D(n2546), .CLK(clk), .Q(
        memoryDataRegister[20]) );
  DFFPOSX1 \ir_reg[20]  ( .D(n1007), .CLK(clk), .Q(N1149) );
  DFFPOSX1 \memoryDataRegister_reg[22]  ( .D(n2550), .CLK(clk), .Q(
        memoryDataRegister[22]) );
  DFFPOSX1 \ir_reg[22]  ( .D(n1006), .CLK(clk), .Q(N1143) );
  DFFPOSX1 \memoryDataRegister_reg[24]  ( .D(n2554), .CLK(clk), .Q(
        memoryDataRegister[24]) );
  DFFPOSX1 \ir_reg[24]  ( .D(n1005), .CLK(clk), .Q(N1137) );
  DFFPOSX1 \memoryDataRegister_reg[26]  ( .D(n2558), .CLK(clk), .Q(
        memoryDataRegister[26]) );
  DFFPOSX1 \ir_reg[26]  ( .D(n1004), .CLK(clk), .Q(N1131) );
  DFFPOSX1 \memoryDataRegister_reg[28]  ( .D(n2562), .CLK(clk), .Q(
        memoryDataRegister[28]) );
  DFFPOSX1 \ir_reg[28]  ( .D(n1003), .CLK(clk), .Q(N1125) );
  DFFPOSX1 \memoryDataRegister_reg[30]  ( .D(n2566), .CLK(clk), .Q(
        memoryDataRegister[30]) );
  DFFPOSX1 \ir_reg[30]  ( .D(n1002), .CLK(clk), .Q(N1119) );
  LATCH \instructionType_tri_enable_reg[2]  ( .CLK(n4358), .D(n2477), .Q(N966)
         );
  LATCH \instructionType_tri_enable_reg[0]  ( .CLK(n4358), .D(n2477), .Q(N972)
         );
  LATCH \instructionType_tri_enable_reg[1]  ( .CLK(n4358), .D(n2477), .Q(N969)
         );
  DFFPOSX1 \memoryDataRegister_reg[1]  ( .D(n2508), .CLK(clk), .Q(
        memoryDataRegister[1]) );
  DFFPOSX1 \ir_reg[1]  ( .D(n1018), .CLK(clk), .Q(N1206) );
  DFFPOSX1 \memoryDataRegister_reg[31]  ( .D(n2504), .CLK(clk), .Q(
        memoryDataRegister[31]) );
  DFFPOSX1 \ir_reg[31]  ( .D(n1033), .CLK(clk), .Q(N1116) );
  LATCH \fpuOperation_reg[1]  ( .CLK(n4359), .D(N721), .Q(fpuOperation[1]) );
  LATCH \fpuOperation_reg[0]  ( .CLK(n4359), .D(N719), .Q(fpuOperation[0]) );
  DFFPOSX1 \aluResultRegister_reg[31]  ( .D(n1850), .CLK(clk), .Q(
        aluResultRegister[31]) );
  DFFPOSX1 \aluResultRegister_reg[0]  ( .D(aluResult[0]), .CLK(clk), .Q(
        aluResultRegister[0]) );
  DFFPOSX1 \aluResultRegister_reg[9]  ( .D(aluResult[9]), .CLK(clk), .Q(
        aluResultRegister[9]) );
  DFFPOSX1 \pc_reg[9]  ( .D(n1467), .CLK(clk), .Q(pc[9]) );
  DFFPOSX1 \aluResultRegister_reg[8]  ( .D(aluResult[8]), .CLK(clk), .Q(
        aluResultRegister[8]) );
  DFFPOSX1 \pc_reg[8]  ( .D(n1466), .CLK(clk), .Q(pc[8]) );
  DFFPOSX1 \aluResultRegister_reg[7]  ( .D(aluResult[7]), .CLK(clk), .Q(
        aluResultRegister[7]) );
  DFFPOSX1 \pc_reg[7]  ( .D(n1465), .CLK(clk), .Q(pc[7]) );
  DFFPOSX1 \aluResultRegister_reg[6]  ( .D(aluResult[6]), .CLK(clk), .Q(
        aluResultRegister[6]) );
  DFFPOSX1 \pc_reg[6]  ( .D(n1464), .CLK(clk), .Q(pc[6]) );
  DFFPOSX1 \aluResultRegister_reg[5]  ( .D(aluResult[5]), .CLK(clk), .Q(
        aluResultRegister[5]) );
  DFFPOSX1 \pc_reg[5]  ( .D(n1463), .CLK(clk), .Q(pc[5]) );
  DFFPOSX1 \aluResultRegister_reg[4]  ( .D(aluResult[4]), .CLK(clk), .Q(
        aluResultRegister[4]) );
  DFFPOSX1 \pc_reg[4]  ( .D(n1462), .CLK(clk), .Q(pc[4]) );
  DFFPOSX1 \aluResultRegister_reg[3]  ( .D(aluResult[3]), .CLK(clk), .Q(
        aluResultRegister[3]) );
  DFFPOSX1 \pc_reg[3]  ( .D(n1461), .CLK(clk), .Q(pc[3]) );
  DFFPOSX1 \aluResultRegister_reg[30]  ( .D(n2225), .CLK(clk), .Q(
        aluResultRegister[30]) );
  DFFPOSX1 \pc_reg[30]  ( .D(n1869), .CLK(clk), .Q(pc[30]) );
  DFFPOSX1 \aluResultRegister_reg[29]  ( .D(aluResult[29]), .CLK(clk), .Q(
        aluResultRegister[29]) );
  DFFPOSX1 \pc_reg[29]  ( .D(n1487), .CLK(clk), .Q(pc[29]) );
  DFFPOSX1 \aluResultRegister_reg[28]  ( .D(aluResult[28]), .CLK(clk), .Q(
        aluResultRegister[28]) );
  DFFPOSX1 \pc_reg[28]  ( .D(n1486), .CLK(clk), .Q(pc[28]) );
  DFFPOSX1 \aluResultRegister_reg[27]  ( .D(aluResult[27]), .CLK(clk), .Q(
        aluResultRegister[27]) );
  DFFPOSX1 \pc_reg[27]  ( .D(n1485), .CLK(clk), .Q(pc[27]) );
  DFFPOSX1 \aluResultRegister_reg[26]  ( .D(aluResult[26]), .CLK(clk), .Q(
        aluResultRegister[26]) );
  DFFPOSX1 \pc_reg[26]  ( .D(n1484), .CLK(clk), .Q(pc[26]) );
  DFFPOSX1 \aluResultRegister_reg[25]  ( .D(aluResult[25]), .CLK(clk), .Q(
        aluResultRegister[25]) );
  DFFPOSX1 \pc_reg[25]  ( .D(n1483), .CLK(clk), .Q(pc[25]) );
  DFFPOSX1 \aluResultRegister_reg[24]  ( .D(aluResult[24]), .CLK(clk), .Q(
        aluResultRegister[24]) );
  DFFPOSX1 \pc_reg[24]  ( .D(n1482), .CLK(clk), .Q(pc[24]) );
  DFFPOSX1 \aluResultRegister_reg[23]  ( .D(aluResult[23]), .CLK(clk), .Q(
        aluResultRegister[23]) );
  DFFPOSX1 \pc_reg[23]  ( .D(n1481), .CLK(clk), .Q(pc[23]) );
  DFFPOSX1 \aluResultRegister_reg[22]  ( .D(aluResult[22]), .CLK(clk), .Q(
        aluResultRegister[22]) );
  DFFPOSX1 \pc_reg[22]  ( .D(n1480), .CLK(clk), .Q(pc[22]) );
  DFFPOSX1 \aluResultRegister_reg[21]  ( .D(aluResult[21]), .CLK(clk), .Q(
        aluResultRegister[21]) );
  DFFPOSX1 \pc_reg[21]  ( .D(n1479), .CLK(clk), .Q(pc[21]) );
  DFFPOSX1 \aluResultRegister_reg[20]  ( .D(aluResult[20]), .CLK(clk), .Q(
        aluResultRegister[20]) );
  DFFPOSX1 \pc_reg[20]  ( .D(n1478), .CLK(clk), .Q(pc[20]) );
  DFFPOSX1 \aluResultRegister_reg[1]  ( .D(aluResult[1]), .CLK(clk), .Q(
        aluResultRegister[1]) );
  DFFPOSX1 \pc_reg[1]  ( .D(n1459), .CLK(clk), .Q(pc[1]) );
  DFFPOSX1 \aluResultRegister_reg[19]  ( .D(aluResult[19]), .CLK(clk), .Q(
        aluResultRegister[19]) );
  DFFPOSX1 \pc_reg[19]  ( .D(n1477), .CLK(clk), .Q(pc[19]) );
  DFFPOSX1 \aluResultRegister_reg[18]  ( .D(aluResult[18]), .CLK(clk), .Q(
        aluResultRegister[18]) );
  DFFPOSX1 \pc_reg[18]  ( .D(n1476), .CLK(clk), .Q(pc[18]) );
  DFFPOSX1 \aluResultRegister_reg[17]  ( .D(aluResult[17]), .CLK(clk), .Q(
        aluResultRegister[17]) );
  DFFPOSX1 \pc_reg[17]  ( .D(n1475), .CLK(clk), .Q(pc[17]) );
  DFFPOSX1 \aluResultRegister_reg[16]  ( .D(aluResult[16]), .CLK(clk), .Q(
        aluResultRegister[16]) );
  DFFPOSX1 \pc_reg[16]  ( .D(n1474), .CLK(clk), .Q(pc[16]) );
  DFFPOSX1 \aluResultRegister_reg[15]  ( .D(aluResult[15]), .CLK(clk), .Q(
        aluResultRegister[15]) );
  DFFPOSX1 \pc_reg[15]  ( .D(n1473), .CLK(clk), .Q(pc[15]) );
  DFFPOSX1 \aluResultRegister_reg[14]  ( .D(aluResult[14]), .CLK(clk), .Q(
        aluResultRegister[14]) );
  DFFPOSX1 \pc_reg[14]  ( .D(n1472), .CLK(clk), .Q(pc[14]) );
  DFFPOSX1 \aluResultRegister_reg[13]  ( .D(aluResult[13]), .CLK(clk), .Q(
        aluResultRegister[13]) );
  DFFPOSX1 \pc_reg[13]  ( .D(n1471), .CLK(clk), .Q(pc[13]) );
  DFFPOSX1 \aluResultRegister_reg[12]  ( .D(aluResult[12]), .CLK(clk), .Q(
        aluResultRegister[12]) );
  DFFPOSX1 \pc_reg[12]  ( .D(n1470), .CLK(clk), .Q(pc[12]) );
  DFFPOSX1 \aluResultRegister_reg[11]  ( .D(aluResult[11]), .CLK(clk), .Q(
        aluResultRegister[11]) );
  DFFPOSX1 \pc_reg[11]  ( .D(n1469), .CLK(clk), .Q(pc[11]) );
  DFFPOSX1 \aluResultRegister_reg[10]  ( .D(aluResult[10]), .CLK(clk), .Q(
        aluResultRegister[10]) );
  DFFPOSX1 \pc_reg[10]  ( .D(n1468), .CLK(clk), .Q(pc[10]) );
  DFFPOSX1 \aluResultRegister_reg[2]  ( .D(aluResult[2]), .CLK(clk), .Q(
        aluResultRegister[2]) );
  DFFPOSX1 \pc_reg[2]  ( .D(n1460), .CLK(clk), .Q(pc[2]) );
  DFFPOSX1 \pc_reg[31]  ( .D(n1870), .CLK(clk), .Q(pc[31]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[16]  ( .A(n2005), .EN(n4031), .Y(
        aluResult[16]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[9]  ( .A(n929), .EN(n4031), .Y(
        aluResult[9]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[7]  ( .A(n925), .EN(n4031), .Y(
        aluResult[7]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[2]  ( .A(n3079), .EN(n4031), .Y(
        aluResult[2]) );
  TBUFX2 \ir_tri[2]  ( .A(n617), .EN(n618), .Y(opcode[2]) );
  TBUFX2 \ir_tri[3]  ( .A(n615), .EN(n616), .Y(opcode[3]) );
  TBUFX2 \ir_tri[4]  ( .A(n613), .EN(n614), .Y(opcode[4]) );
  TBUFX2 \ir_tri[5]  ( .A(n611), .EN(n612), .Y(opcode[5]) );
  TBUFX2 \ir_tri[14]  ( .A(n593), .EN(n594), .Y(funct3[2]) );
  TBUFX2 \aluOperation_tri[3]  ( .A(n3072), .EN(n3561), .Y(aluOperation[3]) );
  OAI21X1 U266 ( .A(funct3[1]), .B(\funct3[0] ), .C(n2220), .Y(n138) );
  AND2X1 U515 ( .A(n4371), .B(n4370), .Y(n217) );
  AOI22X1 U517 ( .A(instructionType[2]), .B(instructionType[1]), .C(n217), .D(
        n4372), .Y(n848) );
  NOR3X1 U904 ( .A(funct7[1]), .B(funct7[0]), .C(n3050), .Y(n978) );
  NAND3X1 U905 ( .A(n978), .B(n1140), .C(n1141), .Y(n977) );
  NAND3X1 U907 ( .A(\funct3[0] ), .B(n1144), .C(n2220), .Y(n980) );
  NAND3X1 U908 ( .A(n3303), .B(n1144), .C(n1138), .Y(n982) );
  NAND3X1 U909 ( .A(funct3[1]), .B(n1145), .C(n1138), .Y(n981) );
  INVX1 U918 ( .A(nextState[4]), .Y(n989) );
  INVX1 U920 ( .A(nextState[0]), .Y(n991) );
  INVX1 U922 ( .A(nextState[3]), .Y(n993) );
  INVX1 U924 ( .A(nextState[2]), .Y(n996) );
  INVX1 U926 ( .A(nextState[1]), .Y(n998) );
  AOI22X1 U1063 ( .A(memoryData[31]), .B(irWrite), .C(n4030), .D(N1116), .Y(
        n1188) );
  AOI22X1 U1064 ( .A(memoryData[30]), .B(irWrite), .C(n4030), .D(N1119), .Y(
        n1190) );
  AOI22X1 U1065 ( .A(memoryData[29]), .B(irWrite), .C(n4030), .D(N1122), .Y(
        n1191) );
  AOI22X1 U1066 ( .A(memoryData[28]), .B(irWrite), .C(n4030), .D(N1125), .Y(
        n1192) );
  AOI22X1 U1067 ( .A(memoryData[27]), .B(irWrite), .C(n4030), .D(N1128), .Y(
        n1193) );
  AOI22X1 U1068 ( .A(memoryData[26]), .B(irWrite), .C(n4030), .D(N1131), .Y(
        n1194) );
  AOI22X1 U1069 ( .A(memoryData[25]), .B(irWrite), .C(n4030), .D(N1134), .Y(
        n1195) );
  AOI22X1 U1070 ( .A(memoryData[24]), .B(irWrite), .C(n4030), .D(N1137), .Y(
        n1196) );
  AOI22X1 U1071 ( .A(memoryData[23]), .B(irWrite), .C(n4030), .D(N1140), .Y(
        n1197) );
  AOI22X1 U1072 ( .A(memoryData[22]), .B(irWrite), .C(n4030), .D(N1143), .Y(
        n1198) );
  AOI22X1 U1073 ( .A(memoryData[21]), .B(irWrite), .C(n4030), .D(N1146), .Y(
        n1199) );
  AOI22X1 U1074 ( .A(memoryData[20]), .B(irWrite), .C(n4030), .D(N1149), .Y(
        n1200) );
  AOI22X1 U1075 ( .A(memoryData[19]), .B(irWrite), .C(n4030), .D(N1152), .Y(
        n1201) );
  AOI22X1 U1076 ( .A(memoryData[18]), .B(irWrite), .C(n4030), .D(N1155), .Y(
        n1202) );
  AOI22X1 U1077 ( .A(memoryData[17]), .B(irWrite), .C(n4030), .D(N1158), .Y(
        n1203) );
  AOI22X1 U1078 ( .A(memoryData[16]), .B(irWrite), .C(n4030), .D(N1161), .Y(
        n1204) );
  AOI22X1 U1079 ( .A(memoryData[15]), .B(irWrite), .C(n4030), .D(N1164), .Y(
        n1205) );
  AOI22X1 U1080 ( .A(memoryData[14]), .B(irWrite), .C(n4030), .D(N1167), .Y(
        n1206) );
  AOI22X1 U1081 ( .A(memoryData[13]), .B(irWrite), .C(n4030), .D(N1170), .Y(
        n1207) );
  AOI22X1 U1082 ( .A(memoryData[12]), .B(irWrite), .C(n4030), .D(N1173), .Y(
        n1208) );
  AOI22X1 U1083 ( .A(memoryData[11]), .B(irWrite), .C(n4030), .D(N1176), .Y(
        n1209) );
  AOI22X1 U1084 ( .A(memoryData[10]), .B(irWrite), .C(n4030), .D(N1179), .Y(
        n1210) );
  AOI22X1 U1085 ( .A(memoryData[9]), .B(irWrite), .C(n4030), .D(N1182), .Y(
        n1211) );
  AOI22X1 U1086 ( .A(memoryData[8]), .B(irWrite), .C(n4030), .D(N1185), .Y(
        n1212) );
  AOI22X1 U1087 ( .A(memoryData[7]), .B(irWrite), .C(n4030), .D(N1188), .Y(
        n1213) );
  AOI22X1 U1204 ( .A(memoryData[5]), .B(irWrite), .C(n4030), .D(N1194), .Y(
        n1275) );
  AOI22X1 U1207 ( .A(memoryData[4]), .B(irWrite), .C(n4030), .D(N1197), .Y(
        n1277) );
  AOI22X1 U1210 ( .A(memoryData[3]), .B(irWrite), .C(n4030), .D(N1200), .Y(
        n1279) );
  AOI22X1 U1213 ( .A(memoryData[2]), .B(irWrite), .C(n4030), .D(N1203), .Y(
        n1281) );
  AOI22X1 U1216 ( .A(memoryData[1]), .B(irWrite), .C(n4030), .D(N1206), .Y(
        n1283) );
  AOI22X1 U1220 ( .A(memoryData[0]), .B(irWrite), .C(n4030), .D(N1209), .Y(
        n1286) );
  AOI22X1 U1221 ( .A(memoryData[6]), .B(irWrite), .C(n4030), .D(N1191), .Y(
        n1287) );
  AOI22X1 U1225 ( .A(RS2[30]), .B(n4029), .C(n4363), .D(memoryDataRegister[30]), .Y(n1288) );
  AOI22X1 U1228 ( .A(RS2[29]), .B(n4029), .C(n4363), .D(memoryDataRegister[29]), .Y(n1293) );
  AOI22X1 U1231 ( .A(RS2[28]), .B(n4029), .C(n4363), .D(memoryDataRegister[28]), .Y(n1295) );
  AOI22X1 U1234 ( .A(RS2[27]), .B(n4029), .C(n4363), .D(memoryDataRegister[27]), .Y(n1297) );
  AOI22X1 U1237 ( .A(RS2[26]), .B(n4029), .C(n4363), .D(memoryDataRegister[26]), .Y(n1299) );
  AOI22X1 U1240 ( .A(RS2[25]), .B(n4029), .C(n4363), .D(memoryDataRegister[25]), .Y(n1301) );
  AOI22X1 U1243 ( .A(RS2[24]), .B(n4029), .C(n4363), .D(memoryDataRegister[24]), .Y(n1303) );
  AOI22X1 U1246 ( .A(RS2[23]), .B(n4029), .C(n4363), .D(memoryDataRegister[23]), .Y(n1305) );
  AOI22X1 U1249 ( .A(RS2[22]), .B(n4029), .C(n4363), .D(memoryDataRegister[22]), .Y(n1307) );
  AOI22X1 U1252 ( .A(RS2[21]), .B(n4029), .C(n4363), .D(memoryDataRegister[21]), .Y(n1309) );
  AOI22X1 U1255 ( .A(RS2[20]), .B(n4029), .C(n4363), .D(memoryDataRegister[20]), .Y(n1311) );
  AOI22X1 U1258 ( .A(RS2[19]), .B(n4029), .C(n4363), .D(memoryDataRegister[19]), .Y(n1313) );
  AOI22X1 U1261 ( .A(RS2[18]), .B(n4029), .C(n4363), .D(memoryDataRegister[18]), .Y(n1315) );
  AOI22X1 U1264 ( .A(RS2[17]), .B(n4029), .C(n4363), .D(memoryDataRegister[17]), .Y(n1317) );
  AOI22X1 U1267 ( .A(RS2[16]), .B(n4029), .C(n4363), .D(memoryDataRegister[16]), .Y(n1319) );
  AOI22X1 U1270 ( .A(RS2[15]), .B(n4029), .C(n4363), .D(memoryDataRegister[15]), .Y(n1321) );
  AOI22X1 U1273 ( .A(RS2[14]), .B(n4029), .C(n4363), .D(memoryDataRegister[14]), .Y(n1323) );
  AOI22X1 U1276 ( .A(RS2[13]), .B(n4029), .C(n4363), .D(memoryDataRegister[13]), .Y(n1325) );
  AOI22X1 U1279 ( .A(RS2[12]), .B(n4029), .C(n4363), .D(memoryDataRegister[12]), .Y(n1327) );
  AOI22X1 U1282 ( .A(RS2[11]), .B(n4029), .C(n4363), .D(memoryDataRegister[11]), .Y(n1329) );
  AOI22X1 U1285 ( .A(RS2[10]), .B(n4029), .C(n4363), .D(memoryDataRegister[10]), .Y(n1331) );
  AOI22X1 U1288 ( .A(RS2[9]), .B(n4029), .C(n4363), .D(memoryDataRegister[9]), 
        .Y(n1333) );
  AOI22X1 U1291 ( .A(RS2[8]), .B(n4029), .C(n4363), .D(memoryDataRegister[8]), 
        .Y(n1335) );
  AOI22X1 U1294 ( .A(RS2[7]), .B(n4029), .C(n4363), .D(memoryDataRegister[7]), 
        .Y(n1337) );
  AOI22X1 U1297 ( .A(RS2[6]), .B(n4029), .C(n4363), .D(memoryDataRegister[6]), 
        .Y(n1339) );
  AOI22X1 U1300 ( .A(RS2[5]), .B(n4029), .C(n4363), .D(memoryDataRegister[5]), 
        .Y(n1341) );
  AOI22X1 U1303 ( .A(RS2[4]), .B(n4029), .C(n4363), .D(memoryDataRegister[4]), 
        .Y(n1343) );
  AOI22X1 U1306 ( .A(RS2[3]), .B(n4029), .C(n4363), .D(memoryDataRegister[3]), 
        .Y(n1345) );
  AOI22X1 U1309 ( .A(RS2[2]), .B(n4029), .C(n4363), .D(memoryDataRegister[2]), 
        .Y(n1347) );
  AOI22X1 U1312 ( .A(RS2[1]), .B(n4029), .C(n4363), .D(memoryDataRegister[1]), 
        .Y(n1349) );
  AOI22X1 U1315 ( .A(RS2[0]), .B(n4029), .C(n4363), .D(memoryDataRegister[0]), 
        .Y(n1351) );
  AOI22X1 U1318 ( .A(RS2[31]), .B(n4029), .C(n4363), .D(memoryDataRegister[31]), .Y(n1353) );
  AOI22X1 U1356 ( .A(instructionOrData), .B(n1156), .C(n1105), .D(n1034), .Y(
        memoryAddress[31]) );
  AOI22X1 U1357 ( .A(instructionOrData), .B(n1157), .C(n1106), .D(n1034), .Y(
        memoryAddress[30]) );
  AOI22X1 U1359 ( .A(instructionOrData), .B(n1158), .C(n1107), .D(n1034), .Y(
        memoryAddress[29]) );
  AOI22X1 U1360 ( .A(instructionOrData), .B(n1159), .C(n1108), .D(n1034), .Y(
        memoryAddress[28]) );
  AOI22X1 U1361 ( .A(instructionOrData), .B(n1160), .C(n1109), .D(n1034), .Y(
        memoryAddress[27]) );
  AOI22X1 U1362 ( .A(instructionOrData), .B(n4038), .C(n1110), .D(n1034), .Y(
        memoryAddress[26]) );
  AOI22X1 U1363 ( .A(instructionOrData), .B(n4040), .C(n1111), .D(n1034), .Y(
        memoryAddress[25]) );
  AOI22X1 U1364 ( .A(instructionOrData), .B(n4042), .C(n1112), .D(n1034), .Y(
        memoryAddress[24]) );
  AOI22X1 U1365 ( .A(instructionOrData), .B(n4044), .C(n1113), .D(n1034), .Y(
        memoryAddress[23]) );
  AOI22X1 U1366 ( .A(instructionOrData), .B(n4046), .C(n1114), .D(n1034), .Y(
        memoryAddress[22]) );
  AOI22X1 U1367 ( .A(instructionOrData), .B(n4048), .C(n1115), .D(n1034), .Y(
        memoryAddress[21]) );
  AOI22X1 U1368 ( .A(instructionOrData), .B(n4050), .C(n1116), .D(n1034), .Y(
        memoryAddress[20]) );
  AOI22X1 U1370 ( .A(instructionOrData), .B(n4052), .C(n1117), .D(n1034), .Y(
        memoryAddress[19]) );
  AOI22X1 U1371 ( .A(instructionOrData), .B(n4054), .C(n1118), .D(n1034), .Y(
        memoryAddress[18]) );
  AOI22X1 U1372 ( .A(instructionOrData), .B(n4056), .C(n1119), .D(n1034), .Y(
        memoryAddress[17]) );
  AOI22X1 U1373 ( .A(instructionOrData), .B(n4058), .C(n1120), .D(n1034), .Y(
        memoryAddress[16]) );
  NOR3X1 U1383 ( .A(aluOperation[2]), .B(aluOperation[3]), .C(n4368), .Y(n1381) );
  NAND3X1 U1425 ( .A(n3530), .B(n3501), .C(n3507), .Y(n1426) );
  NAND3X1 U1426 ( .A(n1430), .B(n4367), .C(n1139), .Y(n1424) );
  AND2X1 U1427 ( .A(n1142), .B(n1143), .Y(n1430) );
  NAND3X1 U1436 ( .A(n2852), .B(n2958), .C(n3037), .Y(n1449) );
  OAI21X1 U1439 ( .A(n1140), .B(n3507), .C(n3530), .Y(N721) );
  OAI21X1 U1441 ( .A(n1141), .B(n3501), .C(n3530), .Y(N719) );
  NAND3X1 U1442 ( .A(funct7[5]), .B(funct7[3]), .C(funct7[2]), .Y(n1427) );
  INVX1 U104 ( .A(funct7[5]), .Y(n1138) );
  INVX1 U110 ( .A(funct3[1]), .Y(n1144) );
  INVX1 U105 ( .A(funct7[4]), .Y(n1139) );
  INVX1 U106 ( .A(funct7[3]), .Y(n1140) );
  INVX1 U107 ( .A(funct7[2]), .Y(n1141) );
  INVX1 U311 ( .A(N1159), .Y(n588) );
  INVX1 U310 ( .A(N1158), .Y(n587) );
  INVX1 U309 ( .A(N1156), .Y(n586) );
  INVX1 U308 ( .A(N1155), .Y(n585) );
  INVX1 U307 ( .A(N1153), .Y(n584) );
  INVX1 U306 ( .A(N1152), .Y(n583) );
  INVX1 U959 ( .A(n1191), .Y(n1032) );
  INVX1 U946 ( .A(n1279), .Y(n1019) );
  INVX1 U948 ( .A(n1213), .Y(n1021) );
  INVX1 U940 ( .A(n1212), .Y(n1013) );
  INVX1 U949 ( .A(n1211), .Y(n1022) );
  INVX1 U939 ( .A(n1210), .Y(n1012) );
  INVX1 U950 ( .A(n1209), .Y(n1023) );
  INVX1 U938 ( .A(n1208), .Y(n1011) );
  INVX1 U951 ( .A(n1207), .Y(n1024) );
  INVX1 U952 ( .A(n1205), .Y(n1025) );
  INVX1 U953 ( .A(n1203), .Y(n1026) );
  INVX1 U954 ( .A(n1201), .Y(n1027) );
  INVX1 U955 ( .A(n1199), .Y(n1028) );
  INVX1 U956 ( .A(n1197), .Y(n1029) );
  INVX1 U957 ( .A(n1195), .Y(n1030) );
  INVX1 U958 ( .A(n1193), .Y(n1031) );
  INVX1 U945 ( .A(n1283), .Y(n1018) );
  INVX1 U944 ( .A(n1286), .Y(n1017) );
  INVX1 U943 ( .A(n1281), .Y(n1016) );
  INVX1 U937 ( .A(n1206), .Y(n1010) );
  INVX1 U941 ( .A(n1287), .Y(n1014) );
  INVX1 U942 ( .A(n1277), .Y(n1015) );
  INVX1 U931 ( .A(n1194), .Y(n1004) );
  INVX1 U930 ( .A(n1192), .Y(n1003) );
  INVX1 U929 ( .A(n1190), .Y(n1002) );
  INVX1 U936 ( .A(n1204), .Y(n1009) );
  INVX1 U960 ( .A(n1188), .Y(n1033) );
  INVX1 U934 ( .A(n1200), .Y(n1007) );
  INVX1 U933 ( .A(n1198), .Y(n1006) );
  INVX1 U932 ( .A(n1196), .Y(n1005) );
  INVX1 U935 ( .A(n1202), .Y(n1008) );
  INVX1 U1031 ( .A(aluResultRegister[31]), .Y(n1156) );
  INVX1 U1032 ( .A(aluResultRegister[30]), .Y(n1157) );
  INVX1 U1033 ( .A(aluResultRegister[29]), .Y(n1158) );
  INVX1 U1034 ( .A(aluResultRegister[28]), .Y(n1159) );
  INVX1 U1035 ( .A(aluResultRegister[27]), .Y(n1160) );
  INVX1 U181 ( .A(memoryReady), .Y(n61) );
  INVX1 U358 ( .A(memoryDataRegister[20]), .Y(n645) );
  INVX1 U354 ( .A(memoryDataRegister[24]), .Y(n637) );
  INVX1 U353 ( .A(memoryDataRegister[25]), .Y(n635) );
  INVX1 U352 ( .A(memoryDataRegister[26]), .Y(n633) );
  INVX1 U351 ( .A(memoryDataRegister[27]), .Y(n631) );
  INVX1 U350 ( .A(memoryDataRegister[28]), .Y(n629) );
  INVX1 U357 ( .A(memoryDataRegister[21]), .Y(n643) );
  INVX1 U348 ( .A(memoryDataRegister[30]), .Y(n625) );
  INVX1 U355 ( .A(memoryDataRegister[23]), .Y(n639) );
  INVX1 U368 ( .A(memoryDataRegister[10]), .Y(n665) );
  INVX1 U367 ( .A(memoryDataRegister[11]), .Y(n663) );
  INVX1 U346 ( .A(memoryDataRegister[31]), .Y(n623) );
  INVX1 U365 ( .A(memoryDataRegister[13]), .Y(n659) );
  INVX1 U364 ( .A(memoryDataRegister[14]), .Y(n657) );
  INVX1 U349 ( .A(memoryDataRegister[29]), .Y(n627) );
  INVX1 U378 ( .A(memoryDataRegister[0]), .Y(n685) );
  INVX1 U361 ( .A(memoryDataRegister[17]), .Y(n651) );
  INVX1 U356 ( .A(memoryDataRegister[22]), .Y(n641) );
  INVX1 U377 ( .A(memoryDataRegister[1]), .Y(n683) );
  INVX1 U376 ( .A(memoryDataRegister[2]), .Y(n681) );
  INVX1 U375 ( .A(memoryDataRegister[3]), .Y(n679) );
  INVX1 U374 ( .A(memoryDataRegister[4]), .Y(n677) );
  INVX1 U373 ( .A(memoryDataRegister[5]), .Y(n675) );
  INVX1 U372 ( .A(memoryDataRegister[6]), .Y(n673) );
  INVX1 U371 ( .A(memoryDataRegister[7]), .Y(n671) );
  INVX1 U370 ( .A(memoryDataRegister[8]), .Y(n669) );
  INVX1 U369 ( .A(memoryDataRegister[9]), .Y(n667) );
  INVX1 U360 ( .A(memoryDataRegister[18]), .Y(n649) );
  INVX1 U359 ( .A(memoryDataRegister[19]), .Y(n647) );
  INVX1 U366 ( .A(memoryDataRegister[12]), .Y(n661) );
  INVX1 U362 ( .A(memoryDataRegister[16]), .Y(n653) );
  INVX1 U363 ( .A(memoryDataRegister[15]), .Y(n655) );
  INVX1 U253 ( .A(N971), .Y(n541) );
  INVX1 U249 ( .A(N965), .Y(n537) );
  INVX1 U251 ( .A(N968), .Y(n539) );
  INVX1 U108 ( .A(funct7[1]), .Y(n1142) );
  INVX1 U109 ( .A(funct7[0]), .Y(n1143) );
  INVX1 U252 ( .A(N969), .Y(n540) );
  INVX1 U250 ( .A(N966), .Y(n538) );
  INVX1 U254 ( .A(N972), .Y(n542) );
  AND2X1 U347 ( .A(memoryReadWrite), .B(memoryEnable), .Y(n624) );
  OR2X2 U1219 ( .A(n4364), .B(irWrite), .Y(n1247) );
  OAI21X1 \sub_x_1100_2/U226  ( .A(n3288), .B(n1825), .C(n3236), .Y(
        \sub_x_1100_2/n170 ) );
  XOR2X1 \sub_x_1100_2/U224  ( .A(n3068), .B(n3656), .Y(
        \arithmetic_logic_unit/N122 ) );
  OAI21X1 \sub_x_1100_2/U219  ( .A(n3529), .B(\sub_x_1100_2/n169 ), .C(n3545), 
        .Y(\sub_x_1100_2/n166 ) );
  OAI21X1 \sub_x_1100_2/U213  ( .A(n3545), .B(n3667), .C(n2229), .Y(
        \sub_x_1100_2/n163 ) );
  AOI21X1 \sub_x_1100_2/U211  ( .A(n2874), .B(\sub_x_1100_2/n170 ), .C(
        \sub_x_1100_2/n163 ), .Y(\sub_x_1100_2/n161 ) );
  XNOR2X1 \sub_x_1100_2/U209  ( .A(\sub_x_1100_2/n166 ), .B(n3118), .Y(
        \arithmetic_logic_unit/N124 ) );
  AOI21X1 \sub_x_1100_2/U202  ( .A(\sub_x_1100_2/n160 ), .B(n3179), .C(n3527), 
        .Y(\sub_x_1100_2/n155 ) );
  OAI21X1 \sub_x_1100_2/U196  ( .A(n3526), .B(n2338), .C(n3233), .Y(
        \sub_x_1100_2/n152 ) );
  AOI21X1 \sub_x_1100_2/U194  ( .A(\sub_x_1100_2/n160 ), .B(n3310), .C(
        \sub_x_1100_2/n152 ), .Y(\sub_x_1100_2/n150 ) );
  XOR2X1 \sub_x_1100_2/U193  ( .A(n3065), .B(n3152), .Y(
        \arithmetic_logic_unit/N126 ) );
  XOR2X1 \sub_x_1100_2/U187  ( .A(n3516), .B(n3150), .Y(
        \arithmetic_logic_unit/N127 ) );
  OAI21X1 \sub_x_1100_2/U182  ( .A(n3669), .B(n3534), .C(n3231), .Y(
        \sub_x_1100_2/n144 ) );
  AOI21X1 \sub_x_1100_2/U180  ( .A(\sub_x_1100_2/n152 ), .B(n3315), .C(
        \sub_x_1100_2/n144 ), .Y(\sub_x_1100_2/n142 ) );
  OAI21X1 \sub_x_1100_2/U165  ( .A(n3542), .B(n2462), .C(n3229), .Y(
        \sub_x_1100_2/n133 ) );
  OAI21X1 \sub_x_1100_2/U161  ( .A(n2451), .B(\sub_x_1100_2/n139 ), .C(
        \sub_x_1100_2/n131 ), .Y(\sub_x_1100_2/n129 ) );
  AOI21X1 \sub_x_1100_2/U153  ( .A(\sub_x_1100_2/n129 ), .B(n3184), .C(n3657), 
        .Y(\sub_x_1100_2/n124 ) );
  OAI21X1 \sub_x_1100_2/U147  ( .A(n3658), .B(n3533), .C(n3227), .Y(
        \sub_x_1100_2/n121 ) );
  AOI21X1 \sub_x_1100_2/U145  ( .A(\sub_x_1100_2/n133 ), .B(n3308), .C(
        \sub_x_1100_2/n121 ), .Y(\sub_x_1100_2/n119 ) );
  OAI21X1 \sub_x_1100_2/U143  ( .A(n3337), .B(\sub_x_1100_2/n139 ), .C(n2459), 
        .Y(\sub_x_1100_2/n117 ) );
  XOR2X1 \sub_x_1100_2/U141  ( .A(n3064), .B(n3148), .Y(
        \arithmetic_logic_unit/N132 ) );
  OAI21X1 \sub_x_1100_2/U128  ( .A(n3524), .B(n3662), .C(n3225), .Y(
        \sub_x_1100_2/n108 ) );
  OAI21X1 \sub_x_1100_2/U124  ( .A(n3163), .B(\sub_x_1100_2/n116 ), .C(
        \sub_x_1100_2/n106 ), .Y(\sub_x_1100_2/n104 ) );
  AOI21X1 \sub_x_1100_2/U116  ( .A(\sub_x_1100_2/n104 ), .B(n2330), .C(n3522), 
        .Y(\sub_x_1100_2/n99 ) );
  OAI21X1 \sub_x_1100_2/U110  ( .A(n3523), .B(n3660), .C(n3223), .Y(
        \sub_x_1100_2/n96 ) );
  AOI21X1 \sub_x_1100_2/U108  ( .A(\sub_x_1100_2/n108 ), .B(n3298), .C(
        \sub_x_1100_2/n96 ), .Y(\sub_x_1100_2/n94 ) );
  OAI21X1 \sub_x_1100_2/U106  ( .A(n3319), .B(n2459), .C(n2686), .Y(
        \sub_x_1100_2/n92 ) );
  AOI21X1 \sub_x_1100_2/U104  ( .A(n2439), .B(n1824), .C(\sub_x_1100_2/n92 ), 
        .Y(\sub_x_1100_2/n90 ) );
  XOR2X1 \sub_x_1100_2/U102  ( .A(n3063), .B(n3146), .Y(
        \arithmetic_logic_unit/N136 ) );
  AOI21X1 \sub_x_1100_2/U95  ( .A(\sub_x_1100_2/n89 ), .B(n3692), .C(n3646), 
        .Y(\sub_x_1100_2/n84 ) );
  AOI21X1 \sub_x_1100_2/U87  ( .A(n2485), .B(n3646), .C(n3639), .Y(
        \sub_x_1100_2/n79 ) );
  OAI21X1 \sub_x_1100_2/U85  ( .A(n2880), .B(n2415), .C(n2685), .Y(
        \sub_x_1100_2/n77 ) );
  XOR2X1 \sub_x_1100_2/U84  ( .A(n3062), .B(n3144), .Y(
        \arithmetic_logic_unit/N138 ) );
  AOI21X1 \sub_x_1100_2/U77  ( .A(\sub_x_1100_2/n77 ), .B(n3687), .C(n3162), 
        .Y(\sub_x_1100_2/n72 ) );
  OAI21X1 \sub_x_1100_2/U71  ( .A(n2414), .B(n3266), .C(n3221), .Y(
        \sub_x_1100_2/n69 ) );
  AOI21X1 \sub_x_1100_2/U63  ( .A(\sub_x_1100_2/n69 ), .B(n3691), .C(n3645), 
        .Y(\sub_x_1100_2/n64 ) );
  XOR2X1 \sub_x_1100_2/U56  ( .A(n3515), .B(n3142), .Y(
        \arithmetic_logic_unit/N142 ) );
  XNOR2X1 \sub_x_1100_2/U48  ( .A(n2213), .B(n3116), .Y(
        \arithmetic_logic_unit/N143 ) );
  XOR2X1 \sub_x_1100_2/U42  ( .A(n2042), .B(n3140), .Y(
        \arithmetic_logic_unit/N144 ) );
  XNOR2X1 \sub_x_1100_2/U34  ( .A(n1815), .B(n3114), .Y(
        \arithmetic_logic_unit/N145 ) );
  XOR2X1 \sub_x_1100_2/U28  ( .A(n3514), .B(n3138), .Y(
        \arithmetic_logic_unit/N146 ) );
  XNOR2X1 \sub_x_1100_2/U20  ( .A(n2214), .B(n3112), .Y(
        \arithmetic_logic_unit/N147 ) );
  XOR2X1 \sub_x_1100_2/U14  ( .A(n2048), .B(n3136), .Y(
        \arithmetic_logic_unit/N148 ) );
  XNOR2X1 \sub_x_1100_2/U6  ( .A(\sub_x_1100_2/n37 ), .B(n3110), .Y(
        \arithmetic_logic_unit/N149 ) );
  FAX1 \sub_x_1100_2/U4  ( .A(n3650), .B(\sub_x_1100_2/A[29] ), .C(
        \sub_x_1100_2/n174 ), .YC(\sub_x_1100_2/n31 ), .YS(
        \arithmetic_logic_unit/N150 ) );
  FAX1 \sub_x_1100_2/U3  ( .A(n3283), .B(\sub_x_1100_2/A[30] ), .C(
        \sub_x_1100_2/n31 ), .YC(\sub_x_1100_2/n30 ), .YS(
        \arithmetic_logic_unit/N151 ) );
  OAI21X1 \add_x_1100_1/U218  ( .A(n2328), .B(n3556), .C(n3212), .Y(
        \add_x_1100_1/n166 ) );
  XOR2X1 \add_x_1100_1/U216  ( .A(n3066), .B(n3557), .Y(
        \arithmetic_logic_unit/N90 ) );
  OAI21X1 \add_x_1100_1/U211  ( .A(n3537), .B(\add_x_1100_1/n165 ), .C(n3541), 
        .Y(\add_x_1100_1/n162 ) );
  OAI21X1 \add_x_1100_1/U205  ( .A(n3541), .B(n2797), .C(n3211), .Y(
        \add_x_1100_1/n159 ) );
  AOI21X1 \add_x_1100_1/U203  ( .A(n2872), .B(\add_x_1100_1/n166 ), .C(
        \add_x_1100_1/n159 ), .Y(\add_x_1100_1/n157 ) );
  XNOR2X1 \add_x_1100_1/U201  ( .A(\add_x_1100_1/n162 ), .B(n3108), .Y(
        \arithmetic_logic_unit/N92 ) );
  AOI21X1 \add_x_1100_1/U194  ( .A(\add_x_1100_1/n156 ), .B(n3177), .C(n3521), 
        .Y(\add_x_1100_1/n151 ) );
  OAI21X1 \add_x_1100_1/U188  ( .A(n3520), .B(n2273), .C(n3208), .Y(
        \add_x_1100_1/n148 ) );
  AOI21X1 \add_x_1100_1/U186  ( .A(\add_x_1100_1/n156 ), .B(n3306), .C(
        \add_x_1100_1/n148 ), .Y(\add_x_1100_1/n146 ) );
  XOR2X1 \add_x_1100_1/U185  ( .A(n3061), .B(n3134), .Y(
        \arithmetic_logic_unit/N94 ) );
  XOR2X1 \add_x_1100_1/U179  ( .A(n3513), .B(n3132), .Y(
        \arithmetic_logic_unit/N95 ) );
  OAI21X1 \add_x_1100_1/U174  ( .A(n2482), .B(n2480), .C(n3206), .Y(
        \add_x_1100_1/n140 ) );
  AOI21X1 \add_x_1100_1/U172  ( .A(\add_x_1100_1/n148 ), .B(n2276), .C(
        \add_x_1100_1/n140 ), .Y(\add_x_1100_1/n138 ) );
  OAI21X1 \add_x_1100_1/U170  ( .A(n2396), .B(n3286), .C(n2684), .Y(
        \add_x_1100_1/n136 ) );
  OAI21X1 \add_x_1100_1/U157  ( .A(n2323), .B(n2463), .C(n3205), .Y(
        \add_x_1100_1/n129 ) );
  OAI21X1 \add_x_1100_1/U153  ( .A(\add_x_1100_1/n126 ), .B(
        \add_x_1100_1/n135 ), .C(\add_x_1100_1/n127 ), .Y(\add_x_1100_1/n125 )
         );
  AOI21X1 \add_x_1100_1/U145  ( .A(\add_x_1100_1/n125 ), .B(
        \add_x_1100_1/n188 ), .C(n3256), .Y(\add_x_1100_1/n120 ) );
  OAI21X1 \add_x_1100_1/U139  ( .A(n3255), .B(n3532), .C(n3203), .Y(
        \add_x_1100_1/n117 ) );
  AOI21X1 \add_x_1100_1/U137  ( .A(\add_x_1100_1/n129 ), .B(n1847), .C(
        \add_x_1100_1/n117 ), .Y(\add_x_1100_1/n115 ) );
  OAI21X1 \add_x_1100_1/U135  ( .A(n2218), .B(\add_x_1100_1/n135 ), .C(n3317), 
        .Y(\add_x_1100_1/n113 ) );
  XOR2X1 \add_x_1100_1/U133  ( .A(n3060), .B(n3130), .Y(
        \arithmetic_logic_unit/N100 ) );
  OAI21X1 \add_x_1100_1/U120  ( .A(n2317), .B(n3664), .C(n3201), .Y(
        \add_x_1100_1/n104 ) );
  OAI21X1 \add_x_1100_1/U116  ( .A(n3175), .B(\add_x_1100_1/n112 ), .C(
        \add_x_1100_1/n102 ), .Y(\add_x_1100_1/n100 ) );
  AOI21X1 \add_x_1100_1/U108  ( .A(\add_x_1100_1/n100 ), .B(\add_x_1100_1/n96 ), .C(n3519), .Y(\add_x_1100_1/n95 ) );
  OAI21X1 \add_x_1100_1/U102  ( .A(n3518), .B(n3531), .C(n3199), .Y(
        \add_x_1100_1/n92 ) );
  AOI21X1 \add_x_1100_1/U100  ( .A(\add_x_1100_1/n104 ), .B(n2287), .C(
        \add_x_1100_1/n92 ), .Y(\add_x_1100_1/n90 ) );
  OAI21X1 \add_x_1100_1/U98  ( .A(n2430), .B(n2457), .C(n2682), .Y(
        \add_x_1100_1/n88 ) );
  AOI21X1 \add_x_1100_1/U96  ( .A(\add_x_1100_1/n136 ), .B(n1857), .C(
        \add_x_1100_1/n88 ), .Y(\add_x_1100_1/n86 ) );
  XOR2X1 \add_x_1100_1/U94  ( .A(n3059), .B(n3128), .Y(
        \arithmetic_logic_unit/N104 ) );
  AOI21X1 \add_x_1100_1/U87  ( .A(\add_x_1100_1/n85 ), .B(n3684), .C(n3161), 
        .Y(\add_x_1100_1/n80 ) );
  AOI21X1 \add_x_1100_1/U79  ( .A(n3683), .B(n3161), .C(n3174), .Y(
        \add_x_1100_1/n75 ) );
  OAI21X1 \add_x_1100_1/U77  ( .A(n2394), .B(n3284), .C(n2681), .Y(
        \add_x_1100_1/n73 ) );
  XOR2X1 \add_x_1100_1/U76  ( .A(n3058), .B(n2434), .Y(
        \arithmetic_logic_unit/N106 ) );
  AOI21X1 \add_x_1100_1/U69  ( .A(n1842), .B(n3682), .C(n3647), .Y(
        \add_x_1100_1/n68 ) );
  OAI21X1 \add_x_1100_1/U63  ( .A(n2423), .B(n2427), .C(n3196), .Y(
        \add_x_1100_1/n65 ) );
  XOR2X1 \add_x_1100_1/U48  ( .A(n3512), .B(n3126), .Y(
        \arithmetic_logic_unit/N110 ) );
  XNOR2X1 \add_x_1100_1/U40  ( .A(n2275), .B(n3636), .Y(
        \arithmetic_logic_unit/N111 ) );
  XOR2X1 \add_x_1100_1/U34  ( .A(n2045), .B(n3124), .Y(
        \arithmetic_logic_unit/N112 ) );
  XNOR2X1 \add_x_1100_1/U26  ( .A(\add_x_1100_1/n49 ), .B(n3638), .Y(
        \arithmetic_logic_unit/N113 ) );
  XOR2X1 \add_x_1100_1/U20  ( .A(n3511), .B(n3122), .Y(
        \arithmetic_logic_unit/N114 ) );
  XNOR2X1 \add_x_1100_1/U12  ( .A(n2224), .B(n3634), .Y(
        \arithmetic_logic_unit/N115 ) );
  XOR2X1 \add_x_1100_1/U6  ( .A(n2050), .B(n3120), .Y(
        \arithmetic_logic_unit/N116 ) );
  FAX1 \add_x_1100_1/U5  ( .A(\lt_x_1100_4/B[28] ), .B(\sub_x_1100_2/A[28] ), 
        .C(\add_x_1100_1/n33 ), .YC(\add_x_1100_1/n32 ), .YS(
        \arithmetic_logic_unit/N117 ) );
  FAX1 \add_x_1100_1/U4  ( .A(\lt_x_1100_4/B[29] ), .B(\sub_x_1100_2/A[29] ), 
        .C(\add_x_1100_1/n32 ), .YC(\add_x_1100_1/n31 ), .YS(
        \arithmetic_logic_unit/N118 ) );
  FAX1 \add_x_1100_1/U3  ( .A(\lt_x_1100_4/B[30] ), .B(\sub_x_1100_2/A[30] ), 
        .C(\add_x_1100_1/n31 ), .YC(\add_x_1100_1/n30 ), .YS(
        \arithmetic_logic_unit/N119 ) );
  TBUFX2 irWrite_tri ( .A(1'b0), .EN(n526), .Y(irWrite) );
  TBUFX2 instructionOrData_tri ( .A(n543), .EN(n544), .Y(instructionOrData) );
  TBUFX2 \instructionType_tri[1]  ( .A(n539), .EN(n540), .Y(instructionType[1]) );
  TBUFX2 \ir_tri[12]  ( .A(n597), .EN(n598), .Y(\funct3[0] ) );
  TBUFX2 \aluOperation_tri[0]  ( .A(n3074), .EN(n3561), .Y(aluOperation[0]) );
  TBUFX2 \memoryData_tri[31]  ( .A(n623), .EN(n624), .Y(memoryData[31]) );
  TBUFX2 \memoryData_tri[30]  ( .A(n625), .EN(n624), .Y(memoryData[30]) );
  TBUFX2 \memoryData_tri[29]  ( .A(n627), .EN(n624), .Y(memoryData[29]) );
  TBUFX2 \memoryData_tri[28]  ( .A(n629), .EN(n624), .Y(memoryData[28]) );
  TBUFX2 \memoryData_tri[27]  ( .A(n631), .EN(n624), .Y(memoryData[27]) );
  TBUFX2 \memoryData_tri[26]  ( .A(n633), .EN(n624), .Y(memoryData[26]) );
  TBUFX2 \memoryData_tri[25]  ( .A(n635), .EN(n624), .Y(memoryData[25]) );
  TBUFX2 \memoryData_tri[24]  ( .A(n637), .EN(n624), .Y(memoryData[24]) );
  TBUFX2 \memoryData_tri[23]  ( .A(n639), .EN(n624), .Y(memoryData[23]) );
  TBUFX2 \memoryData_tri[22]  ( .A(n641), .EN(n624), .Y(memoryData[22]) );
  TBUFX2 \memoryData_tri[21]  ( .A(n643), .EN(n624), .Y(memoryData[21]) );
  TBUFX2 \memoryData_tri[20]  ( .A(n645), .EN(n624), .Y(memoryData[20]) );
  TBUFX2 \memoryData_tri[19]  ( .A(n647), .EN(n624), .Y(memoryData[19]) );
  TBUFX2 \memoryData_tri[18]  ( .A(n649), .EN(n624), .Y(memoryData[18]) );
  TBUFX2 \memoryData_tri[17]  ( .A(n651), .EN(n624), .Y(memoryData[17]) );
  TBUFX2 \memoryData_tri[16]  ( .A(n653), .EN(n624), .Y(memoryData[16]) );
  TBUFX2 \memoryData_tri[15]  ( .A(n655), .EN(n624), .Y(memoryData[15]) );
  TBUFX2 \memoryData_tri[14]  ( .A(n657), .EN(n624), .Y(memoryData[14]) );
  TBUFX2 \memoryData_tri[13]  ( .A(n659), .EN(n624), .Y(memoryData[13]) );
  TBUFX2 \memoryData_tri[12]  ( .A(n661), .EN(n624), .Y(memoryData[12]) );
  TBUFX2 \memoryData_tri[11]  ( .A(n663), .EN(n624), .Y(memoryData[11]) );
  TBUFX2 \memoryData_tri[10]  ( .A(n665), .EN(n624), .Y(memoryData[10]) );
  TBUFX2 \memoryData_tri[9]  ( .A(n667), .EN(n624), .Y(memoryData[9]) );
  TBUFX2 \memoryData_tri[8]  ( .A(n669), .EN(n624), .Y(memoryData[8]) );
  TBUFX2 \memoryData_tri[7]  ( .A(n671), .EN(n624), .Y(memoryData[7]) );
  TBUFX2 \memoryData_tri[6]  ( .A(n673), .EN(n624), .Y(memoryData[6]) );
  TBUFX2 \memoryData_tri[5]  ( .A(n675), .EN(n624), .Y(memoryData[5]) );
  TBUFX2 \memoryData_tri[4]  ( .A(n677), .EN(n624), .Y(memoryData[4]) );
  TBUFX2 \memoryData_tri[3]  ( .A(n679), .EN(n624), .Y(memoryData[3]) );
  TBUFX2 \memoryData_tri[2]  ( .A(n681), .EN(n624), .Y(memoryData[2]) );
  TBUFX2 \memoryData_tri[1]  ( .A(n683), .EN(n624), .Y(memoryData[1]) );
  TBUFX2 \memoryData_tri[0]  ( .A(n685), .EN(n624), .Y(memoryData[0]) );
  TBUFX2 memoryReadWrite_tri ( .A(n517), .EN(n518), .Y(memoryReadWrite) );
  TBUFX2 \arithmetic_logic_unit/result_tri[8]  ( .A(n2003), .EN(n4031), .Y(
        aluResult[8]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[15]  ( .A(n3085), .EN(n4031), .Y(
        aluResult[15]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[23]  ( .A(n3090), .EN(n4031), .Y(
        aluResult[23]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[27]  ( .A(n3093), .EN(n4031), .Y(
        aluResult[27]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[10]  ( .A(n931), .EN(n4031), .Y(
        aluResult[10]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[5]  ( .A(n921), .EN(n4031), .Y(
        aluResult[5]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[0]  ( .A(n2009), .EN(n4031), .Y(
        aluResult[0]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[30]  ( .A(n971), .EN(n4031), .Y(
        aluResult[30]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[4]  ( .A(n2006), .EN(n4031), .Y(
        aluResult[4]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[11]  ( .A(n3082), .EN(n4031), .Y(
        aluResult[11]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[1]  ( .A(n3078), .EN(n4031), .Y(
        aluResult[1]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[17]  ( .A(n3086), .EN(n4031), .Y(
        aluResult[17]) );
  TBUFX2 \instructionType_tri[0]  ( .A(n541), .EN(n542), .Y(instructionType[0]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[12]  ( .A(n2004), .EN(n4031), .Y(
        aluResult[12]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[13]  ( .A(n3084), .EN(n4031), .Y(
        aluResult[13]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[14]  ( .A(n2012), .EN(n4031), .Y(
        aluResult[14]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[18]  ( .A(n947), .EN(n4031), .Y(
        aluResult[18]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[19]  ( .A(n3087), .EN(n4031), .Y(
        aluResult[19]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[20]  ( .A(n2007), .EN(n4031), .Y(
        aluResult[20]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[21]  ( .A(n3089), .EN(n4031), .Y(
        aluResult[21]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[24]  ( .A(n3091), .EN(n4031), .Y(
        aluResult[24]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[25]  ( .A(n3092), .EN(n4031), .Y(
        aluResult[25]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[28]  ( .A(n3094), .EN(n4031), .Y(
        aluResult[28]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[29]  ( .A(n2008), .EN(n4031), .Y(
        aluResult[29]) );
  TBUFX2 \ir_tri[6]  ( .A(n609), .EN(n610), .Y(opcode[6]) );
  TBUFX2 pcWrite_tri ( .A(1'b0), .EN(n524), .Y(pcWrite) );
  TBUFX2 \immediate_generator/immediate_tri[14]  ( .A(n875), .EN(n4032), .Y(
        immediate[14]) );
  TBUFX2 \immediate_generator/immediate_tri[15]  ( .A(n877), .EN(n4032), .Y(
        immediate[15]) );
  TBUFX2 \immediate_generator/immediate_tri[16]  ( .A(n879), .EN(n4032), .Y(
        immediate[16]) );
  TBUFX2 \immediate_generator/immediate_tri[17]  ( .A(n881), .EN(n4032), .Y(
        immediate[17]) );
  TBUFX2 \immediate_generator/immediate_tri[18]  ( .A(n883), .EN(n4032), .Y(
        immediate[18]) );
  TBUFX2 \immediate_generator/immediate_tri[19]  ( .A(n885), .EN(n4032), .Y(
        immediate[19]) );
  TBUFX2 \ir_tri[0]  ( .A(n621), .EN(n622), .Y(\opcode[0] ) );
  TBUFX2 \ir_tri[1]  ( .A(n619), .EN(n620), .Y(\opcode[1] ) );
  TBUFX2 \immediate_generator/immediate_tri[1]  ( .A(n849), .EN(n4032), .Y(
        immediate[1]) );
  TBUFX2 \immediate_generator/immediate_tri[2]  ( .A(n851), .EN(n4032), .Y(
        immediate[2]) );
  TBUFX2 \immediate_generator/immediate_tri[3]  ( .A(n853), .EN(n4032), .Y(
        immediate[3]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[22]  ( .A(n3630), .EN(n4031), .Y(
        aluResult[22]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[26]  ( .A(n3629), .EN(n4031), .Y(
        aluResult[26]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[3]  ( .A(n3080), .EN(n4031), .Y(
        aluResult[3]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[6]  ( .A(n923), .EN(n4031), .Y(
        aluResult[6]) );
  TBUFX2 \ir_tri[13]  ( .A(n595), .EN(n596), .Y(funct3[1]) );
  TBUFX2 \instructionType_tri[2]  ( .A(n537), .EN(n538), .Y(instructionType[2]) );
  TBUFX2 \ir_tri[30]  ( .A(n561), .EN(n562), .Y(funct7[5]) );
  TBUFX2 \ir_tri[25]  ( .A(n571), .EN(n572), .Y(funct7[0]) );
  TBUFX2 \ir_tri[26]  ( .A(n569), .EN(n570), .Y(funct7[1]) );
  TBUFX2 \aluOperation_tri[2]  ( .A(n553), .EN(n3561), .Y(aluOperation[2]) );
  TBUFX2 \ir_tri[27]  ( .A(n567), .EN(n568), .Y(funct7[2]) );
  TBUFX2 \ir_tri[28]  ( .A(n565), .EN(n566), .Y(funct7[3]) );
  TBUFX2 \ir_tri[7]  ( .A(n607), .EN(n608), .Y(ir_7) );
  TBUFX2 \ir_tri[20]  ( .A(n581), .EN(n582), .Y(ir[20]) );
  TBUFX2 \ir_tri[31]  ( .A(n559), .EN(n560), .Y(funct7[6]) );
  TBUFX2 \ir_tri[29]  ( .A(n563), .EN(n564), .Y(funct7[4]) );
  TBUFX2 \aluSrcA_tri[1]  ( .A(n547), .EN(n1845), .Y(aluSrcA[1]) );
  TBUFX2 \ir_tri[21]  ( .A(n579), .EN(n580), .Y(ir[21]) );
  TBUFX2 \ir_tri[22]  ( .A(n577), .EN(n578), .Y(ir[22]) );
  TBUFX2 \ir_tri[23]  ( .A(n575), .EN(n576), .Y(ir[23]) );
  TBUFX2 \ir_tri[24]  ( .A(n573), .EN(n574), .Y(ir[24]) );
  TBUFX2 \aluOperation_tri[1]  ( .A(n3073), .EN(n3561), .Y(aluOperation[1]) );
  TBUFX2 \immediate_generator/immediate_tri[31]  ( .A(n4367), .EN(n4032), .Y(
        immediate[31]) );
  TBUFX2 \immediate_generator/immediate_tri[30]  ( .A(n907), .EN(n4032), .Y(
        immediate[30]) );
  TBUFX2 \immediate_generator/immediate_tri[29]  ( .A(n905), .EN(n4032), .Y(
        immediate[29]) );
  TBUFX2 \immediate_generator/immediate_tri[28]  ( .A(n903), .EN(n4032), .Y(
        immediate[28]) );
  TBUFX2 \immediate_generator/immediate_tri[27]  ( .A(n901), .EN(n4032), .Y(
        immediate[27]) );
  TBUFX2 \immediate_generator/immediate_tri[26]  ( .A(n899), .EN(n4032), .Y(
        immediate[26]) );
  TBUFX2 \immediate_generator/immediate_tri[25]  ( .A(n897), .EN(n4032), .Y(
        immediate[25]) );
  TBUFX2 \immediate_generator/immediate_tri[24]  ( .A(n895), .EN(n4032), .Y(
        immediate[24]) );
  TBUFX2 \immediate_generator/immediate_tri[23]  ( .A(n893), .EN(n4032), .Y(
        immediate[23]) );
  TBUFX2 \immediate_generator/immediate_tri[22]  ( .A(n891), .EN(n4032), .Y(
        immediate[22]) );
  TBUFX2 \immediate_generator/immediate_tri[21]  ( .A(n889), .EN(n4032), .Y(
        immediate[21]) );
  TBUFX2 \immediate_generator/immediate_tri[20]  ( .A(n887), .EN(n4032), .Y(
        immediate[20]) );
  TBUFX2 \immediate_generator/immediate_tri[13]  ( .A(n873), .EN(n4032), .Y(
        immediate[13]) );
  TBUFX2 \immediate_generator/immediate_tri[12]  ( .A(n871), .EN(n4032), .Y(
        immediate[12]) );
  TBUFX2 \immediate_generator/immediate_tri[11]  ( .A(n2473), .EN(n4032), .Y(
        immediate[11]) );
  TBUFX2 \immediate_generator/immediate_tri[10]  ( .A(n3105), .EN(n4032), .Y(
        immediate[10]) );
  TBUFX2 \immediate_generator/immediate_tri[9]  ( .A(n3103), .EN(n4032), .Y(
        immediate[9]) );
  TBUFX2 \immediate_generator/immediate_tri[8]  ( .A(n3101), .EN(n4032), .Y(
        immediate[8]) );
  TBUFX2 \immediate_generator/immediate_tri[7]  ( .A(n3099), .EN(n4032), .Y(
        immediate[7]) );
  TBUFX2 \immediate_generator/immediate_tri[6]  ( .A(n3097), .EN(n4032), .Y(
        immediate[6]) );
  TBUFX2 \immediate_generator/immediate_tri[5]  ( .A(n3095), .EN(n4032), .Y(
        immediate[5]) );
  TBUFX2 \immediate_generator/immediate_tri[4]  ( .A(n855), .EN(n4032), .Y(
        immediate[4]) );
  TBUFX2 \ir_tri[17]  ( .A(n587), .EN(n588), .Y(ir[17]) );
  TBUFX2 \ir_tri[18]  ( .A(n585), .EN(n586), .Y(ir[18]) );
  TBUFX2 \ir_tri[19]  ( .A(n583), .EN(n584), .Y(ir[19]) );
  TBUFX2 \ir_tri[8]  ( .A(n605), .EN(n606), .Y(ir_8) );
  TBUFX2 \ir_tri[9]  ( .A(n603), .EN(n604), .Y(ir_9) );
  TBUFX2 \ir_tri[10]  ( .A(n601), .EN(n602), .Y(ir_10) );
  TBUFX2 \ir_tri[11]  ( .A(n599), .EN(n600), .Y(ir_11) );
  TBUFX2 \ir_tri[15]  ( .A(n591), .EN(n592), .Y(ir[15]) );
  TBUFX2 \ir_tri[16]  ( .A(n589), .EN(n590), .Y(ir[16]) );
  TBUFX2 \immediate_generator/immediate_tri[0]  ( .A(n847), .EN(n4032), .Y(
        immediate[0]) );
  TBUFX2 \nextState_tri[0]  ( .A(n515), .EN(n4362), .Y(nextState[0]) );
  TBUFX2 \nextState_tri[1]  ( .A(n513), .EN(n4362), .Y(nextState[1]) );
  TBUFX2 \nextState_tri[2]  ( .A(n3057), .EN(n4362), .Y(nextState[2]) );
  TBUFX2 \nextState_tri[3]  ( .A(n3055), .EN(n4362), .Y(nextState[3]) );
  TBUFX2 \nextState_tri[4]  ( .A(1'b1), .EN(n4362), .Y(nextState[4]) );
  TBUFX2 \arithmetic_logic_unit/result_tri[31]  ( .A(n2010), .EN(n4031), .Y(
        aluResult[31]) );
  AOI21X1 \sub_x_1100_2/U7  ( .A(\sub_x_1100_2/n37 ), .B(n3686), .C(n3648), 
        .Y(\sub_x_1100_2/n32 ) );
  OAI21X1 \add_x_1100_1/U35  ( .A(n2419), .B(n2046), .C(n3192), .Y(
        \add_x_1100_1/n49 ) );
  OAI21X1 \sub_x_1100_2/U43  ( .A(n2089), .B(n2043), .C(n3217), .Y(
        \sub_x_1100_2/n53 ) );
  TBUFX2 \aluSrcA_tri[0]  ( .A(n3070), .EN(n1845), .Y(aluSrcA[0]) );
  TBUFX2 \aluSrcB_tri[0]  ( .A(n535), .EN(n4361), .Y(aluSrcB[0]) );
  TBUFX2 \aluSrcB_tri[1]  ( .A(n3071), .EN(n4361), .Y(aluSrcB[1]) );
  AOI21X1 U1456 ( .A(\sub_x_1100_2/n53 ), .B(n3689), .C(n3643), .Y(n2058) );
  AOI21X1 U1457 ( .A(n4293), .B(n1557), .C(n1558), .Y(n2005) );
  NAND2X1 U1458 ( .A(n1559), .B(n1560), .Y(n1558) );
  NAND2X1 U1459 ( .A(n2151), .B(n3359), .Y(n1560) );
  AND2X2 U1460 ( .A(n1561), .B(n1562), .Y(n1559) );
  AOI22X1 U1461 ( .A(n1563), .B(n4026), .C(n4027), .D(n1564), .Y(n1562) );
  XNOR2X1 U1462 ( .A(\sub_x_1100_2/n89 ), .B(n1565), .Y(n1564) );
  NAND2X1 U1463 ( .A(n3692), .B(n1566), .Y(n1565) );
  INVX2 U1464 ( .A(n3646), .Y(n1566) );
  XNOR2X1 U1465 ( .A(\add_x_1100_1/n85 ), .B(n1567), .Y(n1563) );
  NAND2X1 U1466 ( .A(n3684), .B(n1568), .Y(n1567) );
  INVX2 U1467 ( .A(n3161), .Y(n1568) );
  AOI21X1 U1468 ( .A(n1569), .B(\lt_x_1100_4/B[16] ), .C(n1570), .Y(n1561) );
  AOI21X1 U1469 ( .A(n2240), .B(n1571), .C(n2084), .Y(n1570) );
  OR2X2 U1470 ( .A(n2241), .B(\lt_x_1100_4/B[16] ), .Y(n1571) );
  NAND2X1 U1471 ( .A(n1572), .B(n2240), .Y(n1569) );
  MUX2X1 U1472 ( .B(n1381), .A(n3704), .S(n2084), .Y(n1572) );
  OAI21X1 U1473 ( .A(n2239), .B(n3338), .C(n1573), .Y(n1557) );
  NAND2X1 U1474 ( .A(n1574), .B(n1575), .Y(n1573) );
  AOI21X1 U1475 ( .A(n3272), .B(n3909), .C(n2236), .Y(n1575) );
  NAND2X1 U1476 ( .A(n3908), .B(n3411), .Y(n1574) );
  AOI21X1 U1477 ( .A(n1576), .B(aluOperation[3]), .C(n1577), .Y(n925) );
  NAND2X1 U1478 ( .A(n1578), .B(n1579), .Y(n1577) );
  AOI21X1 U1479 ( .A(n4026), .B(n1580), .C(n1581), .Y(n1579) );
  NOR2X1 U1480 ( .A(n1582), .B(n3897), .Y(n1581) );
  NAND2X1 U1481 ( .A(n1583), .B(n4293), .Y(n1582) );
  INVX2 U1482 ( .A(n3907), .Y(n1583) );
  XNOR2X1 U1483 ( .A(n1584), .B(n1585), .Y(n1580) );
  OR2X2 U1484 ( .A(n2480), .B(n1586), .Y(n1585) );
  INVX2 U1485 ( .A(n3206), .Y(n1586) );
  OAI21X1 U1486 ( .A(n3536), .B(n3513), .C(n2482), .Y(n1584) );
  AOI21X1 U1487 ( .A(n4027), .B(n1587), .C(n1588), .Y(n1578) );
  NAND2X1 U1488 ( .A(n1589), .B(n1590), .Y(n1588) );
  NAND2X1 U1489 ( .A(n2293), .B(n1591), .Y(n1590) );
  NAND2X1 U1490 ( .A(n1592), .B(n2240), .Y(n1591) );
  MUX2X1 U1491 ( .B(n1381), .A(n3704), .S(n1593), .Y(n1592) );
  INVX2 U1492 ( .A(\sub_x_1100_2/A[7] ), .Y(n1593) );
  NAND2X1 U1493 ( .A(\sub_x_1100_2/A[7] ), .B(n1594), .Y(n1589) );
  NAND2X1 U1494 ( .A(n1595), .B(n2240), .Y(n1594) );
  OR2X2 U1495 ( .A(n2241), .B(n2293), .Y(n1595) );
  XNOR2X1 U1496 ( .A(n1596), .B(n1597), .Y(n1587) );
  NAND2X1 U1497 ( .A(n3231), .B(n1598), .Y(n1597) );
  INVX2 U1498 ( .A(n3534), .Y(n1598) );
  OAI21X1 U1499 ( .A(n3538), .B(n3516), .C(n3669), .Y(n1596) );
  OAI21X1 U1500 ( .A(n2239), .B(n3335), .C(n1599), .Y(n1576) );
  NAND2X1 U1501 ( .A(n1600), .B(n1601), .Y(n1599) );
  NAND2X1 U1502 ( .A(n2286), .B(n3281), .Y(n1601) );
  AOI21X1 U1503 ( .A(n1602), .B(n1603), .C(n1604), .Y(n1600) );
  INVX2 U1504 ( .A(n2239), .Y(n1604) );
  NAND2X1 U1505 ( .A(n2238), .B(n3481), .Y(n1603) );
  AOI21X1 U1506 ( .A(n3500), .B(n2251), .C(n1605), .Y(n1602) );
  INVX2 U1507 ( .A(n3908), .Y(n1605) );
  OAI21X1 U1508 ( .A(n1606), .B(n2052), .C(n1607), .Y(n2049) );
  INVX2 U1509 ( .A(n1608), .Y(n1607) );
  OAI21X1 U1510 ( .A(n3190), .B(n2160), .C(n2161), .Y(n1608) );
  OR2X2 U1511 ( .A(n2160), .B(n2417), .Y(n1606) );
  AOI21X1 U1512 ( .A(n1609), .B(aluOperation[3]), .C(n1610), .Y(n3079) );
  NAND2X1 U1513 ( .A(n1611), .B(n1612), .Y(n1610) );
  NOR2X1 U1514 ( .A(n1613), .B(n1614), .Y(n1612) );
  OAI21X1 U1515 ( .A(n1976), .B(n3342), .C(n1615), .Y(n1614) );
  AOI22X1 U1516 ( .A(n4026), .B(n1616), .C(n1617), .D(n4027), .Y(n1615) );
  XNOR2X1 U1517 ( .A(n1618), .B(\sub_x_1100_2/n169 ), .Y(n1617) );
  NOR2X1 U1518 ( .A(n3544), .B(n3529), .Y(n1618) );
  XOR2X1 U1519 ( .A(\add_x_1100_1/n165 ), .B(n1619), .Y(n1616) );
  NAND2X1 U1520 ( .A(n3541), .B(n2326), .Y(n1619) );
  NOR2X1 U1521 ( .A(n1620), .B(n3651), .Y(n1613) );
  NAND2X1 U1522 ( .A(n1818), .B(n3752), .Y(n1620) );
  NAND2X1 U1523 ( .A(n1621), .B(n1622), .Y(n1611) );
  OAI21X1 U1524 ( .A(n1818), .B(n3651), .C(n1623), .Y(n1622) );
  NAND2X1 U1525 ( .A(n1818), .B(n1381), .Y(n1623) );
  INVX2 U1526 ( .A(n3752), .Y(n1621) );
  OAI21X1 U1527 ( .A(n2239), .B(n3331), .C(n1624), .Y(n1609) );
  NAND2X1 U1528 ( .A(n1625), .B(n1626), .Y(n1624) );
  NAND2X1 U1529 ( .A(n2286), .B(n3468), .Y(n1626) );
  AOI21X1 U1530 ( .A(n1627), .B(n1628), .C(n2236), .Y(n1625) );
  AOI21X1 U1531 ( .A(n1629), .B(n1630), .C(n3909), .Y(n1628) );
  NAND2X1 U1532 ( .A(n3910), .B(n3464), .Y(n1630) );
  AOI21X1 U1533 ( .A(n3462), .B(n1841), .C(n1631), .Y(n1629) );
  INVX2 U1534 ( .A(n2251), .Y(n1631) );
  NAND2X1 U1535 ( .A(n2238), .B(n3499), .Y(n1627) );
  AOI21X1 U1536 ( .A(aluOperation[3]), .B(n1632), .C(n1633), .Y(n931) );
  OAI21X1 U1537 ( .A(n1634), .B(n3326), .C(n1635), .Y(n1633) );
  AOI21X1 U1538 ( .A(\lt_x_1100_4/B[10] ), .B(n1636), .C(n1637), .Y(n1635) );
  NAND2X1 U1539 ( .A(n1638), .B(n1639), .Y(n1637) );
  NAND2X1 U1540 ( .A(\sub_x_1100_2/A[10] ), .B(n1640), .Y(n1639) );
  OAI21X1 U1541 ( .A(\lt_x_1100_4/B[10] ), .B(n2241), .C(n2240), .Y(n1640) );
  AOI22X1 U1542 ( .A(n1641), .B(n4026), .C(n4027), .D(n1642), .Y(n1638) );
  XNOR2X1 U1543 ( .A(\sub_x_1100_2/n129 ), .B(n1643), .Y(n1642) );
  NAND2X1 U1544 ( .A(n3184), .B(n3658), .Y(n1643) );
  XNOR2X1 U1545 ( .A(\add_x_1100_1/n125 ), .B(n1644), .Y(n1641) );
  NAND2X1 U1546 ( .A(n3255), .B(\add_x_1100_1/n188 ), .Y(n1644) );
  NAND2X1 U1547 ( .A(n1645), .B(n2240), .Y(n1636) );
  MUX2X1 U1548 ( .B(n1381), .A(n3704), .S(n1646), .Y(n1645) );
  INVX2 U1549 ( .A(\sub_x_1100_2/A[10] ), .Y(n1646) );
  NAND2X1 U1550 ( .A(n1647), .B(n4293), .Y(n1634) );
  INVX2 U1551 ( .A(n3907), .Y(n1647) );
  NAND2X1 U1552 ( .A(n1648), .B(n1649), .Y(n1632) );
  NAND3X1 U1553 ( .A(n2239), .B(n1650), .C(n1651), .Y(n1649) );
  NAND2X1 U1554 ( .A(n2286), .B(n3275), .Y(n1651) );
  NAND2X1 U1555 ( .A(n3908), .B(n3468), .Y(n1650) );
  OR2X2 U1556 ( .A(n3348), .B(n2239), .Y(n1648) );
  NAND2X1 U1557 ( .A(n3188), .B(n1652), .Y(\add_x_1100_1/n33 ) );
  NAND2X1 U1558 ( .A(n3259), .B(n2049), .Y(n1652) );
  OAI21X1 U1559 ( .A(n1653), .B(n2058), .C(n1654), .Y(n2047) );
  INVX2 U1560 ( .A(n1655), .Y(n1654) );
  OAI21X1 U1561 ( .A(n3215), .B(n2158), .C(n2159), .Y(n1655) );
  OR2X2 U1562 ( .A(n2158), .B(n3261), .Y(n1653) );
  AOI21X1 U1563 ( .A(aluOperation[3]), .B(n1656), .C(n1657), .Y(n929) );
  OAI21X1 U1564 ( .A(n1658), .B(n3330), .C(n1659), .Y(n1657) );
  AOI21X1 U1565 ( .A(\lt_x_1100_4/B[9] ), .B(n1660), .C(n1661), .Y(n1659) );
  NAND2X1 U1566 ( .A(n1662), .B(n1663), .Y(n1661) );
  NAND2X1 U1567 ( .A(n2470), .B(n1664), .Y(n1663) );
  NAND2X1 U1568 ( .A(n1665), .B(n2240), .Y(n1664) );
  OR2X2 U1569 ( .A(n2241), .B(\lt_x_1100_4/B[9] ), .Y(n1665) );
  AOI22X1 U1570 ( .A(n4026), .B(n1666), .C(n4027), .D(n1667), .Y(n1662) );
  XNOR2X1 U1571 ( .A(n1668), .B(n1669), .Y(n1667) );
  NAND2X1 U1572 ( .A(n2461), .B(n3229), .Y(n1669) );
  OAI21X1 U1573 ( .A(n2256), .B(\sub_x_1100_2/n139 ), .C(n3542), .Y(n1668) );
  XNOR2X1 U1574 ( .A(n1670), .B(n1671), .Y(n1666) );
  NAND2X1 U1575 ( .A(n2322), .B(n3205), .Y(n1671) );
  OAI21X1 U1576 ( .A(n2438), .B(\add_x_1100_1/n135 ), .C(n2463), .Y(n1670) );
  NAND2X1 U1577 ( .A(n1672), .B(n2240), .Y(n1660) );
  MUX2X1 U1578 ( .B(n1381), .A(n3704), .S(n1673), .Y(n1672) );
  INVX2 U1579 ( .A(n2469), .Y(n1673) );
  NAND2X1 U1580 ( .A(n1674), .B(n4293), .Y(n1658) );
  INVX2 U1581 ( .A(n3907), .Y(n1674) );
  OAI21X1 U1582 ( .A(n2239), .B(n4014), .C(n1675), .Y(n1656) );
  NAND3X1 U1583 ( .A(n2239), .B(n1676), .C(n1677), .Y(n1675) );
  NAND2X1 U1584 ( .A(n3908), .B(n3495), .Y(n1677) );
  NAND2X1 U1585 ( .A(n2286), .B(n3492), .Y(n1676) );
  NAND2X1 U1586 ( .A(n3213), .B(n1678), .Y(\sub_x_1100_2/n37 ) );
  NAND2X1 U1587 ( .A(n3260), .B(n2047), .Y(n1678) );
  AOI21X1 U1588 ( .A(n4293), .B(n1679), .C(n1680), .Y(n3087) );
  OAI21X1 U1589 ( .A(n1681), .B(n3332), .C(n1682), .Y(n1680) );
  AOI21X1 U1590 ( .A(n1683), .B(n4027), .C(n1684), .Y(n1682) );
  NAND2X1 U1591 ( .A(n1685), .B(n1686), .Y(n1684) );
  NAND2X1 U1592 ( .A(n4026), .B(n1687), .Y(n1686) );
  XOR2X1 U1593 ( .A(n2427), .B(n1688), .Y(n1687) );
  NAND2X1 U1594 ( .A(n3196), .B(n1689), .Y(n1688) );
  INVX2 U1595 ( .A(n2423), .Y(n1689) );
  AOI21X1 U1596 ( .A(n1690), .B(\lt_x_1100_4/B[19] ), .C(n1691), .Y(n1685) );
  NOR2X1 U1597 ( .A(n3759), .B(n1692), .Y(n1691) );
  AOI21X1 U1598 ( .A(n3704), .B(n3247), .C(n3709), .Y(n1692) );
  OAI21X1 U1599 ( .A(n2241), .B(aluOperand1[19]), .C(n1693), .Y(n1690) );
  NOR2X1 U1600 ( .A(n1694), .B(n3709), .Y(n1693) );
  NOR2X1 U1601 ( .A(n1695), .B(n4269), .Y(n1694) );
  INVX2 U1602 ( .A(aluOperand1[19]), .Y(n1695) );
  XOR2X1 U1603 ( .A(n2414), .B(n1696), .Y(n1683) );
  NAND2X1 U1604 ( .A(n3267), .B(n3221), .Y(n1696) );
  OR2X2 U1605 ( .A(n2236), .B(n1697), .Y(n1681) );
  INVX2 U1606 ( .A(aluOperation[3]), .Y(n1697) );
  OAI21X1 U1607 ( .A(n2239), .B(n3344), .C(n1698), .Y(n1679) );
  NAND3X1 U1608 ( .A(n2239), .B(n1699), .C(n1700), .Y(n1698) );
  NAND2X1 U1609 ( .A(n3908), .B(n3420), .Y(n1700) );
  NAND2X1 U1610 ( .A(n3909), .B(n3269), .Y(n1699) );
  AND2X2 U1611 ( .A(n1702), .B(n1701), .Y(n971) );
  NAND2X1 U1612 ( .A(n4026), .B(\arithmetic_logic_unit/N119 ), .Y(n1702) );
  AOI21X1 U1613 ( .A(\arithmetic_logic_unit/N151 ), .B(n4027), .C(n1703), .Y(
        n1701) );
  OAI21X1 U1614 ( .A(n1704), .B(n1705), .C(n1706), .Y(n1703) );
  INVX2 U1615 ( .A(n1707), .Y(n1706) );
  OAI21X1 U1616 ( .A(n1708), .B(n3366), .C(n1709), .Y(n1707) );
  AOI21X1 U1617 ( .A(n1710), .B(\lt_x_1100_4/B[30] ), .C(n1711), .Y(n1709) );
  AOI21X1 U1618 ( .A(n2240), .B(n1712), .C(n1713), .Y(n1711) );
  INVX2 U1619 ( .A(\sub_x_1100_2/A[30] ), .Y(n1713) );
  OR2X2 U1620 ( .A(n2241), .B(\lt_x_1100_4/B[30] ), .Y(n1712) );
  NAND2X1 U1621 ( .A(n1714), .B(n2240), .Y(n1710) );
  AOI21X1 U1622 ( .A(\sub_x_1100_2/A[30] ), .B(n1381), .C(n1715), .Y(n1714) );
  NOR2X1 U1623 ( .A(\sub_x_1100_2/A[30] ), .B(n2241), .Y(n1715) );
  OR2X2 U1624 ( .A(n2236), .B(n2098), .Y(n1708) );
  AOI22X1 U1625 ( .A(n1716), .B(n1717), .C(n3907), .D(n3357), .Y(n1705) );
  NAND2X1 U1626 ( .A(n3909), .B(n3429), .Y(n1717) );
  AOI21X1 U1627 ( .A(n1718), .B(n1719), .C(n2236), .Y(n1716) );
  AOI21X1 U1628 ( .A(n1720), .B(n1721), .C(n3909), .Y(n1719) );
  AOI21X1 U1629 ( .A(n1722), .B(n1723), .C(n2238), .Y(n1721) );
  AOI21X1 U1630 ( .A(\sub_x_1100_2/A[29] ), .B(n1823), .C(n1841), .Y(n1723) );
  NAND2X1 U1631 ( .A(\sub_x_1100_2/A[30] ), .B(n2230), .Y(n1722) );
  NAND2X1 U1632 ( .A(n1841), .B(n3441), .Y(n1720) );
  NAND2X1 U1633 ( .A(n2238), .B(n3438), .Y(n1718) );
  INVX2 U1634 ( .A(n4293), .Y(n1704) );
  NAND2X1 U1635 ( .A(n1725), .B(n1724), .Y(n1869) );
  NAND2X1 U1636 ( .A(n4340), .B(aluResult[30]), .Y(n1725) );
  NAND2X1 U1637 ( .A(pc[30]), .B(n4028), .Y(n1724) );
  AOI21X1 U1638 ( .A(n1726), .B(n1727), .C(n1728), .Y(n2010) );
  NAND2X1 U1639 ( .A(n1729), .B(n1730), .Y(n1728) );
  NAND2X1 U1640 ( .A(n4027), .B(n1731), .Y(n1730) );
  XNOR2X1 U1641 ( .A(\sub_x_1100_2/n30 ), .B(n1732), .Y(n1731) );
  XNOR2X1 U1642 ( .A(\sub_x_1100_2/A[31] ), .B(n3282), .Y(n1732) );
  AOI21X1 U1643 ( .A(n1733), .B(n4293), .C(n1734), .Y(n1729) );
  NAND2X1 U1644 ( .A(n1735), .B(n1736), .Y(n1734) );
  AOI21X1 U1645 ( .A(\sub_x_1100_2/A[31] ), .B(n1737), .C(n1738), .Y(n1736) );
  NOR2X1 U1646 ( .A(n1739), .B(n3368), .Y(n1738) );
  OR2X2 U1647 ( .A(n2236), .B(n2098), .Y(n1739) );
  NAND2X1 U1648 ( .A(n1740), .B(n2240), .Y(n1737) );
  OR2X2 U1649 ( .A(n2241), .B(\lt_x_1100_4/B[31] ), .Y(n1740) );
  NAND2X1 U1650 ( .A(\lt_x_1100_4/B[31] ), .B(n1741), .Y(n1735) );
  NAND2X1 U1651 ( .A(n1742), .B(n2240), .Y(n1741) );
  AOI21X1 U1652 ( .A(\sub_x_1100_2/A[31] ), .B(n1381), .C(n1743), .Y(n1742) );
  NOR2X1 U1653 ( .A(\sub_x_1100_2/A[31] ), .B(n2241), .Y(n1743) );
  NAND2X1 U1654 ( .A(n1744), .B(n1745), .Y(n1733) );
  NAND2X1 U1655 ( .A(n3907), .B(n3358), .Y(n1745) );
  NAND2X1 U1656 ( .A(n1746), .B(n1747), .Y(n1744) );
  NAND2X1 U1657 ( .A(n3909), .B(n3432), .Y(n1747) );
  AOI21X1 U1658 ( .A(n1748), .B(n1749), .C(n2236), .Y(n1746) );
  AOI21X1 U1659 ( .A(n1750), .B(n1751), .C(n2286), .Y(n1749) );
  AOI21X1 U1660 ( .A(n1752), .B(n1753), .C(n2238), .Y(n1751) );
  AND2X2 U1661 ( .A(n1754), .B(n3910), .Y(n1753) );
  NAND2X1 U1662 ( .A(n1823), .B(\sub_x_1100_2/A[30] ), .Y(n1754) );
  NAND2X1 U1663 ( .A(\sub_x_1100_2/A[31] ), .B(n2230), .Y(n1752) );
  NAND2X1 U1664 ( .A(n1841), .B(n3442), .Y(n1750) );
  NAND2X1 U1665 ( .A(n2238), .B(n3440), .Y(n1748) );
  INVX2 U1666 ( .A(n3711), .Y(n1727) );
  XNOR2X1 U1667 ( .A(\add_x_1100_1/n30 ), .B(n1755), .Y(n1726) );
  XNOR2X1 U1668 ( .A(\lt_x_1100_4/B[31] ), .B(\sub_x_1100_2/A[31] ), .Y(n1755)
         );
  AOI21X1 U1669 ( .A(n4026), .B(\arithmetic_logic_unit/N118 ), .C(n1756), .Y(
        n2008) );
  NAND2X1 U1670 ( .A(n1757), .B(n1758), .Y(n1756) );
  NAND2X1 U1671 ( .A(n4027), .B(\arithmetic_logic_unit/N150 ), .Y(n1758) );
  AOI21X1 U1672 ( .A(n1759), .B(n4293), .C(n1760), .Y(n1757) );
  OAI21X1 U1673 ( .A(n1761), .B(n3352), .C(n1762), .Y(n1760) );
  AOI21X1 U1674 ( .A(n1763), .B(\sub_x_1100_2/A[29] ), .C(n1764), .Y(n1762) );
  AOI21X1 U1675 ( .A(n2240), .B(n1765), .C(n3650), .Y(n1764) );
  AOI21X1 U1676 ( .A(\sub_x_1100_2/A[29] ), .B(n1381), .C(n1766), .Y(n1765) );
  NOR2X1 U1677 ( .A(\sub_x_1100_2/A[29] ), .B(n2241), .Y(n1766) );
  NAND2X1 U1678 ( .A(n1767), .B(n2240), .Y(n1763) );
  OR2X2 U1679 ( .A(n2241), .B(\lt_x_1100_4/B[29] ), .Y(n1767) );
  OR2X2 U1680 ( .A(n2236), .B(n2098), .Y(n1761) );
  NAND2X1 U1681 ( .A(n1768), .B(n1769), .Y(n1759) );
  NAND2X1 U1682 ( .A(n3907), .B(n3356), .Y(n1769) );
  NAND2X1 U1683 ( .A(n1770), .B(n1771), .Y(n1768) );
  NAND2X1 U1684 ( .A(n3909), .B(n3426), .Y(n1771) );
  AOI21X1 U1685 ( .A(n1772), .B(n1773), .C(n2236), .Y(n1770) );
  AOI21X1 U1686 ( .A(n1774), .B(n1775), .C(n2286), .Y(n1773) );
  NAND2X1 U1687 ( .A(n3910), .B(n3442), .Y(n1775) );
  AOI21X1 U1688 ( .A(n3439), .B(n1841), .C(n2238), .Y(n1774) );
  NAND2X1 U1689 ( .A(n2238), .B(n3436), .Y(n1772) );
  OR2X1 U1690 ( .A(aluResult[4]), .B(aluResult[1]), .Y(n1799) );
  OR2X1 U1691 ( .A(aluResult[9]), .B(aluResult[7]), .Y(n1795) );
  INVX1 U1692 ( .A(aluResult[19]), .Y(n1798) );
  INVX1 U1693 ( .A(aluResult[12]), .Y(n1797) );
  NOR3X1 U1694 ( .A(aluResult[6]), .B(aluResult[5]), .C(n1799), .Y(n1796) );
  INVX1 U1695 ( .A(aluResult[13]), .Y(n1792) );
  INVX1 U1696 ( .A(aluResult[18]), .Y(n1791) );
  NOR3X1 U1697 ( .A(aluResult[2]), .B(aluResult[3]), .C(aluResult[8]), .Y(
        n1790) );
  NOR3X1 U1698 ( .A(aluResult[16]), .B(aluResult[10]), .C(n1795), .Y(n1794) );
  NAND3X1 U1699 ( .A(n1796), .B(n1797), .C(n1798), .Y(n1793) );
  NAND3X1 U1700 ( .A(n1790), .B(n1791), .C(n1792), .Y(n1789) );
  OR2X1 U1701 ( .A(aluResult[20]), .B(aluResult[14]), .Y(n1808) );
  INVX1 U1702 ( .A(n1794), .Y(n1801) );
  INVX1 U1703 ( .A(n1793), .Y(n1803) );
  BUFX2 U1704 ( .A(n1789), .Y(n1807) );
  OR2X1 U1705 ( .A(aluResult[11]), .B(aluResult[17]), .Y(n1788) );
  OR2X1 U1706 ( .A(n1801), .B(n1808), .Y(n1809) );
  INVX1 U1707 ( .A(n1803), .Y(n1804) );
  INVX1 U1708 ( .A(aluResult[21]), .Y(n1787) );
  NOR3X1 U1709 ( .A(n1788), .B(n1807), .C(aluResult[15]), .Y(n1786) );
  NOR3X1 U1710 ( .A(aluResult[0]), .B(n1804), .C(n1809), .Y(n1785) );
  NAND3X1 U1711 ( .A(n1785), .B(n1786), .C(n1787), .Y(n1784) );
  BUFX2 U1712 ( .A(n1784), .Y(n1806) );
  INVX1 U1713 ( .A(aluResult[25]), .Y(n1783) );
  INVX1 U1714 ( .A(aluResult[24]), .Y(n1782) );
  NOR3X1 U1715 ( .A(aluResult[22]), .B(n1806), .C(aluResult[23]), .Y(n1781) );
  NAND3X1 U1716 ( .A(n1781), .B(n1782), .C(n1783), .Y(n1780) );
  BUFX2 U1717 ( .A(n1780), .Y(n1805) );
  INVX2 U1718 ( .A(aluResult[29]), .Y(n1779) );
  INVX2 U1719 ( .A(aluResult[28]), .Y(n1778) );
  NOR3X1 U1720 ( .A(aluResult[26]), .B(n1805), .C(aluResult[27]), .Y(n1777) );
  NAND3X1 U1721 ( .A(n1777), .B(n1778), .C(n1779), .Y(n1776) );
  BUFX2 U1722 ( .A(n1776), .Y(n1802) );
  INVX1 U1723 ( .A(n2211), .Y(n1800) );
  NOR3X1 U1724 ( .A(n1800), .B(n1802), .C(n2225), .Y(n1554) );
  NAND2X1 U1725 ( .A(n1811), .B(n1810), .Y(n1870) );
  NAND2X1 U1726 ( .A(n4340), .B(aluResult[31]), .Y(n1811) );
  NAND2X1 U1727 ( .A(pc[31]), .B(n4028), .Y(n1810) );
  AND2X2 U1728 ( .A(n3663), .B(n2315), .Y(n1812) );
  INVX2 U1729 ( .A(n1812), .Y(n3175) );
  INVX4 U1730 ( .A(n3663), .Y(n3664) );
  INVX2 U1731 ( .A(n3693), .Y(n2266) );
  INVX4 U1732 ( .A(n3693), .Y(n1813) );
  OAI21X1 U1733 ( .A(n2882), .B(n3287), .C(n2687), .Y(n1814) );
  BUFX2 U1734 ( .A(\sub_x_1100_2/n53 ), .Y(n1815) );
  OAI21X1 U1735 ( .A(n2880), .B(n2415), .C(n2685), .Y(n1816) );
  INVX4 U1736 ( .A(n2278), .Y(n3693) );
  INVX1 U1737 ( .A(n3693), .Y(n1833) );
  INVX1 U1738 ( .A(n3693), .Y(n1832) );
  INVX2 U1739 ( .A(n2280), .Y(n2243) );
  INVX4 U1740 ( .A(n2350), .Y(n2280) );
  INVX1 U1741 ( .A(\ashr_1100_6/SH[2] ), .Y(n1817) );
  INVX2 U1742 ( .A(n1817), .Y(n1818) );
  INVX4 U1743 ( .A(n3707), .Y(\ashr_1100_6/SH[2] ) );
  INVX2 U1744 ( .A(n3749), .Y(n1819) );
  INVX2 U1745 ( .A(n3763), .Y(n1820) );
  BUFX2 U1746 ( .A(aluOperand1[13]), .Y(\sub_x_1100_2/A[13] ) );
  INVX1 U1747 ( .A(n3712), .Y(n1821) );
  BUFX2 U1748 ( .A(n3287), .Y(n1822) );
  BUFX2 U1749 ( .A(\ashr_1100_6/SH[0] ), .Y(n1823) );
  AND2X2 U1750 ( .A(n2280), .B(RS2[1]), .Y(n2374) );
  AND2X2 U1751 ( .A(n3320), .B(n2333), .Y(n1824) );
  INVX2 U1752 ( .A(n2350), .Y(n2216) );
  INVX2 U1753 ( .A(n2350), .Y(n2215) );
  INVX2 U1754 ( .A(n2280), .Y(n2283) );
  INVX4 U1755 ( .A(\lt_x_1100_4/B[13] ), .Y(n2264) );
  INVX2 U1756 ( .A(n3655), .Y(n1825) );
  BUFX2 U1757 ( .A(n2329), .Y(n1826) );
  BUFX2 U1758 ( .A(n2262), .Y(n1827) );
  INVX1 U1759 ( .A(\lt_x_1100_4/B[15] ), .Y(n2262) );
  INVX4 U1760 ( .A(n2349), .Y(n3562) );
  INVX1 U1761 ( .A(n2363), .Y(n1828) );
  BUFX2 U1762 ( .A(N1174), .Y(n1829) );
  BUFX2 U1763 ( .A(aluSrcB[0]), .Y(n1830) );
  INVX2 U1764 ( .A(n2261), .Y(n1831) );
  AND2X2 U1765 ( .A(n4030), .B(n1829), .Y(n3603) );
  INVX4 U1766 ( .A(\lt_x_1100_4/B[9] ), .Y(n2260) );
  INVX2 U1767 ( .A(n4089), .Y(n3694) );
  INVX2 U1768 ( .A(N1200), .Y(n615) );
  BUFX2 U1769 ( .A(n4115), .Y(n1834) );
  INVX2 U1770 ( .A(n2243), .Y(n2282) );
  OR2X2 U1771 ( .A(\sub_x_1100_2/A[8] ), .B(\lt_x_1100_4/B[8] ), .Y(n3535) );
  INVX1 U1772 ( .A(n3673), .Y(n3674) );
  INVX1 U1773 ( .A(n3559), .Y(n3558) );
  OR2X1 U1774 ( .A(n2796), .B(n2219), .Y(n3056) );
  OR2X1 U1775 ( .A(n2115), .B(n1941), .Y(n2011) );
  AND2X1 U1776 ( .A(n1862), .B(n1879), .Y(n1940) );
  AND2X1 U1777 ( .A(n1863), .B(n2127), .Y(n3084) );
  AND2X1 U1778 ( .A(n2222), .B(n3171), .Y(n2488) );
  AND2X1 U1779 ( .A(n2223), .B(n4323), .Y(n2489) );
  AND2X1 U1780 ( .A(n2239), .B(n1871), .Y(n1988) );
  OR2X1 U1781 ( .A(n3342), .B(n2239), .Y(n2099) );
  AND2X1 U1782 ( .A(n4293), .B(n2239), .Y(n2130) );
  INVX2 U1783 ( .A(n2286), .Y(n3908) );
  AND2X1 U1784 ( .A(n2212), .B(n4365), .Y(n2921) );
  INVX1 U1785 ( .A(n3713), .Y(n4023) );
  INVX1 U1786 ( .A(n3714), .Y(n4029) );
  BUFX2 U1787 ( .A(\ashr_1100_6/SH[1] ), .Y(n1841) );
  INVX1 U1788 ( .A(n4293), .Y(n2100) );
  INVX1 U1789 ( .A(aluOperand1[20]), .Y(n2154) );
  INVX1 U1790 ( .A(aluOperand1[16]), .Y(n2084) );
  INVX1 U1791 ( .A(n2230), .Y(n2226) );
  INVX1 U1792 ( .A(n2390), .Y(n2298) );
  AND2X1 U1793 ( .A(\sub_x_1100_2/A[0] ), .B(n2193), .Y(n2192) );
  AND2X1 U1794 ( .A(n3704), .B(n1856), .Y(n2080) );
  INVX1 U1795 ( .A(n3250), .Y(n3249) );
  AND2X1 U1796 ( .A(n2251), .B(n1889), .Y(n2170) );
  AND2X1 U1797 ( .A(n2900), .B(n3910), .Y(n2171) );
  AND2X1 U1798 ( .A(n3282), .B(\sub_x_1100_2/A[31] ), .Y(n2179) );
  INVX1 U1799 ( .A(\sub_x_1100_2/A[8] ), .Y(n2069) );
  INVX1 U1800 ( .A(n2191), .Y(n2190) );
  INVX1 U1801 ( .A(n3688), .Y(n2158) );
  INVX1 U1802 ( .A(n3681), .Y(n2160) );
  INVX1 U1803 ( .A(aluResultRegister[9]), .Y(n1855) );
  AND2X1 U1804 ( .A(n3766), .B(n1895), .Y(n2183) );
  INVX1 U1805 ( .A(n3690), .Y(n2087) );
  INVX1 U1806 ( .A(n3679), .Y(n2142) );
  INVX1 U1807 ( .A(n3251), .Y(\lt_x_1100_4/B[12] ) );
  INVX1 U1808 ( .A(n3162), .Y(n2096) );
  INVX1 U1809 ( .A(n3647), .Y(n2097) );
  AND2X1 U1810 ( .A(n4104), .B(aluOperation[0]), .Y(n2172) );
  INVX1 U1811 ( .A(opcode[4]), .Y(n4147) );
  INVX1 U1812 ( .A(n3160), .Y(n2148) );
  AND2X1 U1813 ( .A(n3239), .B(n2183), .Y(n2181) );
  AND2X1 U1814 ( .A(n3239), .B(n2183), .Y(n2200) );
  AND2X1 U1815 ( .A(n2078), .B(n2079), .Y(n2077) );
  OR2X1 U1816 ( .A(n1939), .B(n3790), .Y(n2039) );
  INVX1 U1817 ( .A(n2313), .Y(n3531) );
  INVX1 U1818 ( .A(n3645), .Y(n2150) );
  INVX1 U1819 ( .A(n3184), .Y(n3183) );
  AND2X1 U1820 ( .A(n1860), .B(n2108), .Y(n1946) );
  INVX1 U1821 ( .A(n1856), .Y(n1846) );
  INVX1 U1822 ( .A(opcode[3]), .Y(n1848) );
  AND2X1 U1823 ( .A(n2829), .B(n2206), .Y(n2205) );
  AND2X1 U1824 ( .A(n2924), .B(n2247), .Y(n2182) );
  AND2X1 U1825 ( .A(n2189), .B(n1893), .Y(n2187) );
  AND2X1 U1826 ( .A(n3325), .B(n2231), .Y(n2206) );
  AND2X1 U1827 ( .A(n1868), .B(n2182), .Y(n1950) );
  AND2X1 U1828 ( .A(n2167), .B(n1927), .Y(n1886) );
  AND2X1 U1829 ( .A(n1864), .B(n1883), .Y(n1948) );
  AND2X1 U1830 ( .A(n2187), .B(n1891), .Y(n1952) );
  AND2X1 U1831 ( .A(n1861), .B(n1875), .Y(n1959) );
  INVX1 U1832 ( .A(n3169), .Y(n2177) );
  INVX1 U1833 ( .A(n3170), .Y(n2197) );
  INVX1 U1834 ( .A(n2246), .Y(n2203) );
  INVX1 U1835 ( .A(n2249), .Y(n2207) );
  OR2X1 U1836 ( .A(n2212), .B(n61), .Y(n4122) );
  MUX2X1 U1837 ( .B(n1381), .A(n3704), .S(n3760), .Y(n1835) );
  AND2X1 U1838 ( .A(n2240), .B(n1835), .Y(n1920) );
  INVX1 U1839 ( .A(n4322), .Y(n1836) );
  NOR3X1 U1840 ( .A(n2309), .B(n3558), .C(n1836), .Y(n4358) );
  INVX1 U1841 ( .A(n3716), .Y(n4030) );
  AOI22X1 U1842 ( .A(immediate[18]), .B(n2306), .C(RS2[18]), .D(n2281), .Y(
        n1837) );
  INVX1 U1843 ( .A(n1837), .Y(\lt_x_1100_4/B[18] ) );
  AOI22X1 U1844 ( .A(aluResult[16]), .B(n4340), .C(pc[16]), .D(n4028), .Y(
        n1838) );
  INVX1 U1845 ( .A(n1838), .Y(n1474) );
  AOI22X1 U1846 ( .A(aluResult[28]), .B(n4340), .C(pc[28]), .D(n4028), .Y(
        n1839) );
  INVX1 U1847 ( .A(n1839), .Y(n1486) );
  AOI22X1 U1848 ( .A(aluResult[8]), .B(n4340), .C(pc[8]), .D(n4028), .Y(n1840)
         );
  INVX1 U1849 ( .A(n1840), .Y(n1466) );
  INVX2 U1850 ( .A(n3705), .Y(\ashr_1100_6/SH[1] ) );
  OAI21X1 U1851 ( .A(n2394), .B(n2428), .C(n2681), .Y(n1842) );
  BUFX2 U1852 ( .A(n4361), .Y(n1843) );
  BUFX2 U1853 ( .A(n4332), .Y(n1844) );
  NOR3X1 U1854 ( .A(n2360), .B(n2367), .C(n2288), .Y(n1845) );
  OR2X2 U1855 ( .A(n3660), .B(n2250), .Y(n3297) );
  INVX1 U1856 ( .A(\lt_x_1100_4/B[12] ), .Y(n1856) );
  INVX2 U1857 ( .A(n2390), .Y(n2302) );
  INVX1 U1858 ( .A(n2319), .Y(n1847) );
  INVX1 U1859 ( .A(n1848), .Y(n1849) );
  INVX2 U1860 ( .A(n2211), .Y(n1850) );
  AND2X1 U1861 ( .A(n4102), .B(immediate[2]), .Y(n2643) );
  INVX4 U1862 ( .A(n2435), .Y(n2437) );
  AND2X2 U1863 ( .A(n2412), .B(n2272), .Y(n1851) );
  INVX2 U1864 ( .A(n2272), .Y(n3720) );
  AND2X2 U1865 ( .A(n2262), .B(n2060), .Y(n3224) );
  INVX2 U1866 ( .A(n4036), .Y(n1854) );
  INVX1 U1867 ( .A(aluSrcA[1]), .Y(n1852) );
  OAI21X1 U1868 ( .A(n1854), .B(n1855), .C(n4071), .Y(n1853) );
  INVX1 U1869 ( .A(n4102), .Y(n4025) );
  INVX1 U1870 ( .A(\sub_x_1100_2/A[14] ), .Y(n2120) );
  AND2X2 U1871 ( .A(n2318), .B(n2429), .Y(n1857) );
  AND2X1 U1872 ( .A(n4102), .B(immediate[0]), .Y(n2646) );
  INVX4 U1873 ( .A(n3252), .Y(\lt_x_1100_4/B[11] ) );
  BUFX2 U1874 ( .A(n2261), .Y(n1858) );
  AND2X1 U1875 ( .A(n4102), .B(immediate[1]), .Y(n2644) );
  INVX2 U1876 ( .A(n2309), .Y(n3548) );
  OR2X1 U1877 ( .A(n4334), .B(n2269), .Y(n2361) );
  INVX2 U1878 ( .A(n2361), .Y(n2362) );
  OR2X2 U1879 ( .A(n3726), .B(n3724), .Y(n3673) );
  INVX1 U1880 ( .A(aluOperation[3]), .Y(n2098) );
  INVX1 U1881 ( .A(n3711), .Y(n4026) );
  INVX2 U1882 ( .A(n3710), .Y(n4027) );
  INVX2 U1883 ( .A(n3655), .Y(n3656) );
  OR2X2 U1884 ( .A(n2060), .B(n2262), .Y(n3659) );
  INVX1 U1885 ( .A(n2461), .Y(n2462) );
  INVX1 U1886 ( .A(n2334), .Y(n3533) );
  OR2X2 U1887 ( .A(\sub_x_1100_2/A[11] ), .B(n3252), .Y(n2334) );
  INVX1 U1888 ( .A(n3641), .Y(n2159) );
  INVX1 U1889 ( .A(n3156), .Y(n2161) );
  INVX1 U1890 ( .A(n3159), .Y(n2143) );
  INVX1 U1891 ( .A(n3642), .Y(n2088) );
  INVX1 U1892 ( .A(n3200), .Y(n3201) );
  INVX2 U1893 ( .A(n3671), .Y(n2290) );
  BUFX4 U1894 ( .A(aluOperand1[11]), .Y(\sub_x_1100_2/A[11] ) );
  OR2X1 U1895 ( .A(n3709), .B(n2112), .Y(n2106) );
  INVX1 U1896 ( .A(n2179), .Y(n2199) );
  AND2X2 U1897 ( .A(n3672), .B(n3720), .Y(n2355) );
  BUFX2 U1898 ( .A(n2064), .Y(n1859) );
  BUFX2 U1899 ( .A(n2107), .Y(n1860) );
  BUFX2 U1900 ( .A(n2101), .Y(n1861) );
  BUFX2 U1901 ( .A(n2116), .Y(n1862) );
  BUFX2 U1902 ( .A(n2126), .Y(n1863) );
  BUFX2 U1903 ( .A(n2131), .Y(n1864) );
  AND2X2 U1904 ( .A(\lt_x_1100_4/B[18] ), .B(n1921), .Y(n1865) );
  INVX1 U1905 ( .A(n1865), .Y(n1866) );
  AND2X1 U1906 ( .A(n3740), .B(n3239), .Y(n1867) );
  INVX1 U1907 ( .A(n1867), .Y(n1868) );
  BUFX2 U1908 ( .A(n2114), .Y(n1871) );
  AND2X2 U1909 ( .A(\sub_x_1100_2/A[8] ), .B(n2065), .Y(n1872) );
  INVX1 U1910 ( .A(n1872), .Y(n1873) );
  AND2X1 U1911 ( .A(n3908), .B(n3417), .Y(n1874) );
  INVX1 U1912 ( .A(n1874), .Y(n1875) );
  AND2X2 U1913 ( .A(aluOperand1[18]), .B(n2102), .Y(n1876) );
  INVX1 U1914 ( .A(n1876), .Y(n1877) );
  AND2X2 U1915 ( .A(n2130), .B(n3357), .Y(n1878) );
  INVX1 U1916 ( .A(n1878), .Y(n1879) );
  AND2X1 U1917 ( .A(n2236), .B(n3366), .Y(n1880) );
  INVX1 U1918 ( .A(n1880), .Y(n1881) );
  AND2X1 U1919 ( .A(n4027), .B(n2132), .Y(n1882) );
  INVX1 U1920 ( .A(n1882), .Y(n1883) );
  AND2X2 U1921 ( .A(n2331), .B(\sub_x_1100_2/n117 ), .Y(n1884) );
  INVX1 U1922 ( .A(n1884), .Y(n1885) );
  INVX1 U1923 ( .A(n1886), .Y(n1887) );
  AND2X1 U1924 ( .A(n2171), .B(n1931), .Y(n1888) );
  INVX1 U1925 ( .A(n1888), .Y(n1889) );
  AND2X1 U1926 ( .A(n2188), .B(n4027), .Y(n1890) );
  INVX1 U1927 ( .A(n1890), .Y(n1891) );
  AND2X1 U1928 ( .A(n2190), .B(n4026), .Y(n1892) );
  INVX1 U1929 ( .A(n1892), .Y(n1893) );
  AND2X2 U1930 ( .A(aluOperand1[16]), .B(n2263), .Y(n1894) );
  INVX1 U1931 ( .A(n1894), .Y(n1895) );
  BUFX2 U1932 ( .A(n2093), .Y(n1896) );
  BUFX2 U1933 ( .A(n2063), .Y(n1897) );
  BUFX2 U1934 ( .A(n2073), .Y(n1898) );
  BUFX2 U1935 ( .A(n2105), .Y(n1899) );
  BUFX2 U1936 ( .A(n2175), .Y(n1900) );
  BUFX2 U1937 ( .A(n2178), .Y(n1901) );
  BUFX2 U1938 ( .A(n2186), .Y(n1902) );
  BUFX2 U1939 ( .A(n2195), .Y(n1903) );
  BUFX2 U1940 ( .A(n2198), .Y(n1904) );
  AND2X1 U1941 ( .A(n1932), .B(n1919), .Y(n1905) );
  INVX1 U1942 ( .A(n1905), .Y(n1906) );
  AND2X1 U1943 ( .A(n1937), .B(n1917), .Y(n1907) );
  INVX1 U1944 ( .A(n1907), .Y(n1908) );
  AND2X1 U1945 ( .A(n2236), .B(n3362), .Y(n1909) );
  INVX1 U1946 ( .A(n1909), .Y(n1910) );
  AND2X1 U1947 ( .A(n4027), .B(n2124), .Y(n1911) );
  INVX1 U1948 ( .A(n1911), .Y(n1912) );
  AND2X1 U1949 ( .A(n1933), .B(n1923), .Y(n1913) );
  INVX1 U1950 ( .A(n1913), .Y(n1914) );
  AND2X1 U1951 ( .A(n1934), .B(n1925), .Y(n1915) );
  INVX1 U1952 ( .A(n1915), .Y(n1916) );
  BUFX2 U1953 ( .A(n2083), .Y(n1917) );
  AND2X1 U1954 ( .A(n3908), .B(n3460), .Y(n1918) );
  INVX1 U1955 ( .A(n1918), .Y(n1919) );
  INVX1 U1956 ( .A(n1920), .Y(n1921) );
  AND2X1 U1957 ( .A(n2286), .B(n3279), .Y(n1922) );
  INVX1 U1958 ( .A(n1922), .Y(n1923) );
  AND2X1 U1959 ( .A(n3908), .B(n3423), .Y(n1924) );
  INVX1 U1960 ( .A(n1924), .Y(n1925) );
  AND2X1 U1961 ( .A(n1935), .B(n1929), .Y(n1926) );
  INVX1 U1962 ( .A(n1926), .Y(n1927) );
  AND2X1 U1963 ( .A(n2286), .B(n3460), .Y(n1928) );
  INVX1 U1964 ( .A(n1928), .Y(n1929) );
  AND2X1 U1965 ( .A(n3722), .B(n4022), .Y(n1930) );
  INVX1 U1966 ( .A(n1930), .Y(n1931) );
  BUFX2 U1967 ( .A(n2070), .Y(n1932) );
  BUFX2 U1968 ( .A(n2129), .Y(n1933) );
  BUFX2 U1969 ( .A(n2157), .Y(n1934) );
  BUFX2 U1970 ( .A(n2168), .Y(n1935) );
  AND2X1 U1971 ( .A(n3908), .B(n3484), .Y(n1936) );
  INVX1 U1972 ( .A(n1936), .Y(n1937) );
  AND2X1 U1973 ( .A(n2252), .B(n2235), .Y(n1938) );
  INVX1 U1974 ( .A(n1938), .Y(n1939) );
  INVX1 U1975 ( .A(n1940), .Y(n1941) );
  BUFX2 U1976 ( .A(n2145), .Y(n1942) );
  BUFX2 U1977 ( .A(n2164), .Y(n1943) );
  AND2X2 U1978 ( .A(n1859), .B(n1873), .Y(n1944) );
  INVX1 U1979 ( .A(n1944), .Y(n1945) );
  INVX1 U1980 ( .A(n1946), .Y(n1947) );
  INVX1 U1981 ( .A(n1948), .Y(n1949) );
  INVX1 U1982 ( .A(n1950), .Y(n1951) );
  INVX1 U1983 ( .A(n1952), .Y(n1953) );
  BUFX2 U1984 ( .A(n2146), .Y(n1954) );
  BUFX2 U1985 ( .A(n2165), .Y(n1955) );
  BUFX2 U1986 ( .A(n2169), .Y(n1956) );
  AND2X1 U1987 ( .A(n2068), .B(n2240), .Y(n1957) );
  INVX1 U1988 ( .A(n1957), .Y(n1958) );
  INVX1 U1989 ( .A(n1959), .Y(n1960) );
  AND2X1 U1990 ( .A(n2208), .B(n2747), .Y(n1961) );
  INVX1 U1991 ( .A(n1961), .Y(n1962) );
  AND2X1 U1992 ( .A(n1841), .B(n3464), .Y(n1963) );
  INVX1 U1993 ( .A(n1963), .Y(n1964) );
  AND2X1 U1994 ( .A(n2238), .B(n3463), .Y(n1965) );
  INVX1 U1995 ( .A(n1965), .Y(n1966) );
  AND2X1 U1996 ( .A(n2870), .B(n2858), .Y(n1967) );
  INVX1 U1997 ( .A(n1967), .Y(n1968) );
  BUFX2 U1998 ( .A(n2119), .Y(n1969) );
  BUFX2 U1999 ( .A(n2123), .Y(n1970) );
  BUFX2 U2000 ( .A(n2135), .Y(n1971) );
  BUFX2 U2001 ( .A(n2153), .Y(n1972) );
  AND2X1 U2002 ( .A(n2040), .B(n3379), .Y(n1973) );
  INVX1 U2003 ( .A(n1973), .Y(n1974) );
  AND2X1 U2004 ( .A(n2239), .B(n4293), .Y(n1975) );
  INVX1 U2005 ( .A(n1975), .Y(n1976) );
  AND2X1 U2006 ( .A(n2040), .B(n3380), .Y(n1977) );
  INVX1 U2007 ( .A(n1977), .Y(n1978) );
  AND2X1 U2008 ( .A(n2238), .B(n3459), .Y(n1979) );
  INVX1 U2009 ( .A(n1979), .Y(n1980) );
  AND2X1 U2010 ( .A(n4027), .B(n2149), .Y(n1981) );
  INVX1 U2011 ( .A(n1981), .Y(n1982) );
  AND2X1 U2012 ( .A(n2172), .B(n2173), .Y(n1983) );
  INVX1 U2013 ( .A(n1983), .Y(n1984) );
  BUFX2 U2014 ( .A(n2174), .Y(n1985) );
  BUFX2 U2015 ( .A(n2194), .Y(n1986) );
  BUFX2 U2016 ( .A(n2204), .Y(n1987) );
  INVX1 U2017 ( .A(n1988), .Y(n1989) );
  AND2X2 U2018 ( .A(aluOperation[3]), .B(n1881), .Y(n1990) );
  INVX1 U2019 ( .A(n1990), .Y(n1991) );
  BUFX2 U2020 ( .A(n2201), .Y(n1992) );
  AND2X1 U2021 ( .A(n2251), .B(n3463), .Y(n1993) );
  INVX1 U2022 ( .A(n1993), .Y(n1994) );
  AND2X1 U2023 ( .A(n4026), .B(n2147), .Y(n1995) );
  INVX1 U2024 ( .A(n1995), .Y(n1996) );
  AND2X2 U2025 ( .A(n1866), .B(n1877), .Y(n1997) );
  INVX1 U2026 ( .A(n1997), .Y(n1998) );
  BUFX2 U2027 ( .A(n2090), .Y(n1999) );
  BUFX2 U2028 ( .A(n1104), .Y(n3725) );
  BUFX2 U2029 ( .A(n2138), .Y(n2000) );
  AND2X2 U2030 ( .A(n3524), .B(n1885), .Y(n2001) );
  INVX1 U2031 ( .A(n2001), .Y(n2002) );
  BUFX2 U2032 ( .A(n927), .Y(n2003) );
  BUFX2 U2033 ( .A(n3083), .Y(n2004) );
  BUFX2 U2034 ( .A(n3081), .Y(n2006) );
  BUFX2 U2035 ( .A(n3088), .Y(n2007) );
  BUFX2 U2036 ( .A(n3107), .Y(n2009) );
  INVX1 U2037 ( .A(n2011), .Y(n2012) );
  OR2X2 U2038 ( .A(n2256), .B(n3543), .Y(n2013) );
  INVX1 U2039 ( .A(n2013), .Y(n2014) );
  OR2X2 U2040 ( .A(n2438), .B(n2324), .Y(n2015) );
  INVX1 U2041 ( .A(n2015), .Y(n2016) );
  AND2X2 U2042 ( .A(n2317), .B(\add_x_1100_1/n186 ), .Y(n2017) );
  INVX1 U2043 ( .A(n2017), .Y(n2018) );
  AND2X1 U2044 ( .A(n3687), .B(n2096), .Y(n2019) );
  INVX1 U2045 ( .A(n2019), .Y(n2020) );
  AND2X1 U2046 ( .A(n3682), .B(n2097), .Y(n2021) );
  INVX1 U2047 ( .A(n2021), .Y(n2022) );
  AND2X2 U2048 ( .A(n3520), .B(n3177), .Y(n2023) );
  INVX1 U2049 ( .A(n2023), .Y(n2024) );
  AND2X2 U2050 ( .A(n3179), .B(n3526), .Y(n2025) );
  INVX1 U2051 ( .A(n2025), .Y(n2026) );
  AND2X2 U2052 ( .A(\add_x_1100_1/n96 ), .B(n3518), .Y(n2027) );
  INVX1 U2053 ( .A(n2027), .Y(n2028) );
  AND2X2 U2054 ( .A(n3523), .B(n2330), .Y(n2029) );
  INVX1 U2055 ( .A(n2029), .Y(n2030) );
  AND2X2 U2056 ( .A(n3225), .B(n3661), .Y(n2031) );
  INVX1 U2057 ( .A(n2031), .Y(n2032) );
  OR2X2 U2058 ( .A(n3664), .B(n3200), .Y(n2033) );
  INVX1 U2059 ( .A(n2033), .Y(n2034) );
  AND2X1 U2060 ( .A(n3680), .B(n2148), .Y(n2035) );
  INVX1 U2061 ( .A(n2035), .Y(n2036) );
  AND2X1 U2062 ( .A(n3691), .B(n2150), .Y(n2037) );
  INVX1 U2063 ( .A(n2037), .Y(n2038) );
  INVX1 U2064 ( .A(n2039), .Y(n2040) );
  OR2X2 U2065 ( .A(n2086), .B(n2085), .Y(n2041) );
  INVX1 U2066 ( .A(n2041), .Y(n2042) );
  INVX1 U2067 ( .A(n2041), .Y(n2043) );
  OR2X2 U2068 ( .A(n2141), .B(n2140), .Y(n2044) );
  INVX1 U2069 ( .A(n2044), .Y(n2045) );
  INVX1 U2070 ( .A(n2044), .Y(n2046) );
  INVX1 U2071 ( .A(n2047), .Y(n2048) );
  INVX1 U2072 ( .A(n2049), .Y(n2050) );
  BUFX2 U2073 ( .A(n2426), .Y(n2051) );
  BUFX2 U2074 ( .A(n2425), .Y(n2052) );
  AND2X1 U2075 ( .A(\lt_x_1100_4/B[31] ), .B(n3751), .Y(n2053) );
  INVX1 U2076 ( .A(n2053), .Y(n2054) );
  OR2X1 U2077 ( .A(\sub_x_1100_2/A[30] ), .B(n3283), .Y(n2055) );
  INVX1 U2078 ( .A(n2055), .Y(n2056) );
  BUFX2 U2079 ( .A(n2180), .Y(n2057) );
  BUFX2 U2080 ( .A(\sub_x_1100_2/n64 ), .Y(n2059) );
  BUFX2 U2081 ( .A(aluOperand1[15]), .Y(n2060) );
  AND2X2 U2082 ( .A(n3252), .B(\sub_x_1100_2/A[11] ), .Y(n3228) );
  BUFX4 U2083 ( .A(aluOperand1[7]), .Y(\sub_x_1100_2/A[7] ) );
  INVX2 U2084 ( .A(n2359), .Y(n2360) );
  AOI21X1 U2085 ( .A(aluOperation[3]), .B(n2061), .C(n2062), .Y(n927) );
  OAI21X1 U2086 ( .A(n1976), .B(n3329), .C(n1897), .Y(n2062) );
  AOI21X1 U2087 ( .A(\lt_x_1100_4/B[8] ), .B(n1958), .C(n1945), .Y(n2063) );
  OAI21X1 U2088 ( .A(\lt_x_1100_4/B[8] ), .B(n2241), .C(n2240), .Y(n2065) );
  AOI22X1 U2089 ( .A(n4026), .B(n2066), .C(n4027), .D(n2067), .Y(n2064) );
  XNOR2X1 U2090 ( .A(\sub_x_1100_2/n139 ), .B(n2014), .Y(n2067) );
  XNOR2X1 U2091 ( .A(\add_x_1100_1/n135 ), .B(n2016), .Y(n2066) );
  MUX2X1 U2092 ( .B(n1381), .A(n3704), .S(n2069), .Y(n2068) );
  OAI21X1 U2093 ( .A(n2239), .B(n4011), .C(n1906), .Y(n2061) );
  AOI21X1 U2094 ( .A(n3453), .B(n2286), .C(n2236), .Y(n2070) );
  AOI21X1 U2095 ( .A(aluOperation[3]), .B(n2071), .C(n2072), .Y(n3083) );
  OAI21X1 U2096 ( .A(n1976), .B(n3328), .C(n1898), .Y(n2072) );
  AOI21X1 U2097 ( .A(n2074), .B(n4027), .C(n2075), .Y(n2073) );
  OAI21X1 U2098 ( .A(n3711), .B(n2076), .C(n2077), .Y(n2075) );
  OAI21X1 U2099 ( .A(n2080), .B(n3709), .C(\sub_x_1100_2/A[12] ), .Y(n2079) );
  OAI21X1 U2100 ( .A(n3709), .B(n2081), .C(n1846), .Y(n2078) );
  MUX2X1 U2101 ( .B(n2241), .A(n4269), .S(\sub_x_1100_2/A[12] ), .Y(n2081) );
  XNOR2X1 U2102 ( .A(\add_x_1100_1/n112 ), .B(n2018), .Y(n2076) );
  XNOR2X1 U2103 ( .A(\sub_x_1100_2/n116 ), .B(n2082), .Y(n2074) );
  AND2X2 U2104 ( .A(n2331), .B(n3524), .Y(n2082) );
  OAI21X1 U2105 ( .A(n2239), .B(n3336), .C(n1908), .Y(n2071) );
  AOI21X1 U2106 ( .A(n3483), .B(n2286), .C(n2236), .Y(n2083) );
  NOR3X1 U2107 ( .A(n3264), .B(n2087), .C(n2059), .Y(n2086) );
  OAI21X1 U2108 ( .A(n3219), .B(n2087), .C(n2088), .Y(n2085) );
  INVX1 U2109 ( .A(n3263), .Y(n2089) );
  NOR3X1 U2110 ( .A(n1998), .B(n1999), .C(n2091), .Y(n947) );
  OAI21X1 U2111 ( .A(n2092), .B(n3331), .C(n1896), .Y(n2091) );
  AOI22X1 U2112 ( .A(n4026), .B(n2094), .C(n4027), .D(n2095), .Y(n2093) );
  XNOR2X1 U2113 ( .A(n1816), .B(n2020), .Y(n2095) );
  XNOR2X1 U2114 ( .A(\add_x_1100_1/n73 ), .B(n2022), .Y(n2094) );
  OR2X2 U2115 ( .A(n2236), .B(n2098), .Y(n2092) );
  AOI21X1 U2116 ( .A(n2099), .B(n1960), .C(n2100), .Y(n2090) );
  AOI21X1 U2117 ( .A(n3268), .B(n3909), .C(n2236), .Y(n2101) );
  OAI21X1 U2118 ( .A(\lt_x_1100_4/B[18] ), .B(n2241), .C(n2240), .Y(n2102) );
  AOI21X1 U2119 ( .A(\add_x_1100_1/n65 ), .B(n3680), .C(n3160), .Y(n2426) );
  AOI21X1 U2120 ( .A(aluOperation[3]), .B(n2103), .C(n2104), .Y(n3081) );
  OAI21X1 U2121 ( .A(n1976), .B(n3347), .C(n1899), .Y(n2104) );
  AOI21X1 U2122 ( .A(n2106), .B(n2236), .C(n1947), .Y(n2105) );
  OAI21X1 U2123 ( .A(n2109), .B(n3709), .C(\sub_x_1100_2/A[4] ), .Y(n2108) );
  AND2X2 U2124 ( .A(n3704), .B(n3670), .Y(n2109) );
  AOI22X1 U2125 ( .A(n4027), .B(n2110), .C(n4026), .D(n2111), .Y(n2107) );
  XNOR2X1 U2126 ( .A(\add_x_1100_1/n156 ), .B(n2024), .Y(n2111) );
  XNOR2X1 U2127 ( .A(\sub_x_1100_2/n160 ), .B(n2026), .Y(n2110) );
  MUX2X1 U2128 ( .B(n2241), .A(n4269), .S(\sub_x_1100_2/A[4] ), .Y(n2112) );
  OAI21X1 U2129 ( .A(n2113), .B(n1989), .C(n1910), .Y(n2103) );
  NAND3X1 U2130 ( .A(n3908), .B(n1980), .C(n1994), .Y(n2114) );
  AND2X2 U2131 ( .A(n3484), .B(n2286), .Y(n2113) );
  AOI21X1 U2132 ( .A(n2117), .B(n4026), .C(n2118), .Y(n2116) );
  OAI21X1 U2133 ( .A(n1969), .B(n2120), .C(n2121), .Y(n2118) );
  OAI21X1 U2134 ( .A(n3709), .B(n2122), .C(n3249), .Y(n2121) );
  MUX2X1 U2135 ( .B(n2241), .A(n4269), .S(\sub_x_1100_2/A[14] ), .Y(n2122) );
  AOI21X1 U2136 ( .A(n3704), .B(n3250), .C(n3709), .Y(n2119) );
  XNOR2X1 U2137 ( .A(\add_x_1100_1/n100 ), .B(n2028), .Y(n2117) );
  OAI21X1 U2138 ( .A(n1970), .B(n1991), .C(n1912), .Y(n2115) );
  XNOR2X1 U2139 ( .A(\sub_x_1100_2/n104 ), .B(n2030), .Y(n2124) );
  AOI21X1 U2140 ( .A(n2286), .B(n3490), .C(n2125), .Y(n2123) );
  OAI21X1 U2141 ( .A(n3909), .B(n3280), .C(n2239), .Y(n2125) );
  OAI21X1 U2142 ( .A(n2239), .B(n3352), .C(n1914), .Y(n2128) );
  AOI21X1 U2143 ( .A(n3489), .B(n3908), .C(n2236), .Y(n2129) );
  AOI21X1 U2144 ( .A(n3356), .B(n2130), .C(n1949), .Y(n2126) );
  XNOR2X1 U2145 ( .A(n2002), .B(n2032), .Y(n2132) );
  AOI21X1 U2146 ( .A(n2133), .B(n4026), .C(n2134), .Y(n2131) );
  OAI21X1 U2147 ( .A(n1971), .B(n3763), .C(n2136), .Y(n2134) );
  OAI21X1 U2148 ( .A(n3709), .B(n2137), .C(\lt_x_1100_4/B[13] ), .Y(n2136) );
  MUX2X1 U2149 ( .B(n2241), .A(n4269), .S(n1820), .Y(n2137) );
  AOI21X1 U2150 ( .A(n3704), .B(n2264), .C(n3709), .Y(n2135) );
  XNOR2X1 U2151 ( .A(n2000), .B(n2034), .Y(n2133) );
  AOI21X1 U2152 ( .A(\add_x_1100_1/n113 ), .B(\add_x_1100_1/n186 ), .C(n2316), 
        .Y(n2138) );
  AND2X2 U2153 ( .A(aluOperation[3]), .B(n2128), .Y(n2139) );
  INVX1 U2154 ( .A(n2139), .Y(n2127) );
  NOR3X1 U2155 ( .A(n2421), .B(n2142), .C(n2051), .Y(n2141) );
  OAI21X1 U2156 ( .A(n3194), .B(n2142), .C(n2143), .Y(n2140) );
  AOI21X1 U2157 ( .A(n2144), .B(n4293), .C(n1942), .Y(n3088) );
  NAND3X1 U2158 ( .A(n1954), .B(n1982), .C(n1996), .Y(n2145) );
  XNOR2X1 U2159 ( .A(\add_x_1100_1/n65 ), .B(n2036), .Y(n2147) );
  XNOR2X1 U2160 ( .A(\sub_x_1100_2/n69 ), .B(n2038), .Y(n2149) );
  AOI21X1 U2161 ( .A(n3362), .B(n2151), .C(n2152), .Y(n2146) );
  OAI21X1 U2162 ( .A(n1972), .B(n2154), .C(n2155), .Y(n2152) );
  OAI21X1 U2163 ( .A(n3709), .B(n2156), .C(\lt_x_1100_4/B[20] ), .Y(n2155) );
  MUX2X1 U2164 ( .B(n2241), .A(n4269), .S(aluOperand1[20]), .Y(n2156) );
  AOI21X1 U2165 ( .A(n3704), .B(n3246), .C(n3709), .Y(n2153) );
  AND2X2 U2166 ( .A(n2239), .B(aluOperation[3]), .Y(n2151) );
  OAI21X1 U2167 ( .A(n2239), .B(n3347), .C(n1916), .Y(n2144) );
  AOI21X1 U2168 ( .A(n3271), .B(n3909), .C(n2236), .Y(n2157) );
  AOI21X1 U2169 ( .A(\add_x_1100_1/n49 ), .B(n3678), .C(n3158), .Y(n2425) );
  INVX1 U2170 ( .A(\sub_x_1100_2/n32 ), .Y(\sub_x_1100_2/n174 ) );
  AOI21X1 U2171 ( .A(n2162), .B(n2163), .C(n1943), .Y(n3107) );
  NAND3X1 U2172 ( .A(n1955), .B(n1984), .C(n2166), .Y(n2164) );
  AOI21X1 U2173 ( .A(n1966), .B(n1956), .C(n2236), .Y(n2168) );
  AOI21X1 U2174 ( .A(n1964), .B(n2170), .C(n3909), .Y(n2169) );
  OAI21X1 U2175 ( .A(n1974), .B(n1985), .C(n1900), .Y(n2173) );
  AOI21X1 U2176 ( .A(n3379), .B(n3794), .C(n2176), .Y(n2175) );
  OAI21X1 U2177 ( .A(n2177), .B(n2877), .C(n1901), .Y(n2176) );
  AOI21X1 U2178 ( .A(n2054), .B(n2056), .C(n2179), .Y(n2178) );
  AOI21X1 U2179 ( .A(n2057), .B(n2181), .C(n1951), .Y(n2174) );
  AOI21X1 U2180 ( .A(n2184), .B(\sub_x_1100_2/A[0] ), .C(n2185), .Y(n2165) );
  OAI21X1 U2181 ( .A(n1976), .B(n3338), .C(n1902), .Y(n2185) );
  AOI21X1 U2182 ( .A(n3709), .B(n4022), .C(n1953), .Y(n2186) );
  XNOR2X1 U2183 ( .A(\sub_x_1100_2/A[0] ), .B(n2230), .Y(n2188) );
  OAI21X1 U2184 ( .A(n4022), .B(\sub_x_1100_2/A[0] ), .C(n3557), .Y(n2191) );
  OAI21X1 U2185 ( .A(n2192), .B(n3656), .C(n3704), .Y(n2189) );
  INVX2 U2186 ( .A(n1823), .Y(n2193) );
  OAI21X1 U2187 ( .A(n4269), .B(n2193), .C(n2240), .Y(n2184) );
  OAI21X1 U2188 ( .A(n1978), .B(n1986), .C(n1903), .Y(n2163) );
  AOI21X1 U2189 ( .A(n3380), .B(n3794), .C(n2196), .Y(n2195) );
  OAI21X1 U2190 ( .A(n2197), .B(n2877), .C(n1904), .Y(n2196) );
  AOI21X1 U2191 ( .A(n2056), .B(n2199), .C(n2053), .Y(n2198) );
  AOI21X1 U2192 ( .A(n2057), .B(n2200), .C(n1951), .Y(n2194) );
  AOI22X1 U2193 ( .A(n2257), .B(aluOperand1[17]), .C(n1992), .D(n2202), .Y(
        n2180) );
  OAI21X1 U2194 ( .A(n2203), .B(n1987), .C(n2205), .Y(n2202) );
  AOI21X1 U2195 ( .A(n2746), .B(n1962), .C(n2207), .Y(n2204) );
  OAI21X1 U2196 ( .A(n2878), .B(n3771), .C(n2650), .Y(n2208) );
  AOI21X1 U2197 ( .A(n1968), .B(n3312), .C(n3735), .Y(n2201) );
  NOR3X1 U2198 ( .A(n4368), .B(aluOperation[0]), .C(n4369), .Y(n2162) );
  OR2X1 U2199 ( .A(n2239), .B(n2209), .Y(n2167) );
  AND2X2 U2200 ( .A(aluOperation[3]), .B(n1887), .Y(n2210) );
  INVX1 U2201 ( .A(n2210), .Y(n2166) );
  INVX1 U2202 ( .A(n3359), .Y(n2209) );
  INVX2 U2203 ( .A(aluResult[31]), .Y(n2211) );
  OR2X2 U2204 ( .A(n4322), .B(n3725), .Y(n4131) );
  OR2X2 U2205 ( .A(n3725), .B(n3724), .Y(n2466) );
  OR2X2 U2206 ( .A(n3725), .B(n4366), .Y(n2309) );
  BUFX2 U2207 ( .A(n3675), .Y(n2212) );
  OAI21X1 U2208 ( .A(n3264), .B(n2059), .C(n3219), .Y(n2213) );
  OAI21X1 U2209 ( .A(n3261), .B(n2058), .C(n3215), .Y(n2214) );
  BUFX2 U2210 ( .A(n1814), .Y(n2217) );
  INVX2 U2211 ( .A(n2366), .Y(n2367) );
  INVX1 U2212 ( .A(\lt_x_1100_4/B[5] ), .Y(n2261) );
  AND2X2 U2213 ( .A(\sub_x_1100_2/n227 ), .B(\sub_x_1100_2/A[7] ), .Y(n3232)
         );
  AND2X2 U2214 ( .A(n2264), .B(\sub_x_1100_2/A[13] ), .Y(n3226) );
  OR2X2 U2215 ( .A(\sub_x_1100_2/A[13] ), .B(n2264), .Y(n3661) );
  AND2X2 U2216 ( .A(\lt_x_1100_4/B[13] ), .B(aluOperand1[13]), .Y(n3200) );
  OR2X2 U2217 ( .A(aluOperand1[13]), .B(\lt_x_1100_4/B[13] ), .Y(n3663) );
  AND2X2 U2218 ( .A(\lt_x_1100_4/B[15] ), .B(n2060), .Y(n3198) );
  INVX1 U2219 ( .A(n2318), .Y(n2218) );
  BUFX2 U2220 ( .A(n2360), .Y(n2219) );
  BUFX2 U2221 ( .A(funct3[2]), .Y(n2220) );
  BUFX2 U2222 ( .A(n4147), .Y(n2221) );
  BUFX2 U2223 ( .A(opcode[4]), .Y(n2222) );
  OR2X2 U2224 ( .A(n3533), .B(n3183), .Y(n3307) );
  BUFX2 U2225 ( .A(n1849), .Y(n2223) );
  OAI21X1 U2226 ( .A(n2417), .B(n3511), .C(n3190), .Y(n2224) );
  OR2X2 U2227 ( .A(n3172), .B(n3546), .Y(n2450) );
  BUFX2 U2228 ( .A(n1821), .Y(n2286) );
  INVX2 U2229 ( .A(n3256), .Y(n3255) );
  INVX4 U2230 ( .A(n3657), .Y(n3658) );
  AND2X2 U2231 ( .A(n2233), .B(aluOperand1[10]), .Y(n3657) );
  OR2X2 U2232 ( .A(n2233), .B(aluOperand1[10]), .Y(n3184) );
  AND2X2 U2233 ( .A(n2257), .B(aluOperand1[17]), .Y(n3639) );
  AND2X2 U2234 ( .A(\lt_x_1100_4/B[17] ), .B(aluOperand1[17]), .Y(n3174) );
  AND2X2 U2235 ( .A(n2263), .B(aluOperand1[16]), .Y(n3646) );
  AND2X2 U2236 ( .A(\lt_x_1100_4/B[16] ), .B(aluOperand1[16]), .Y(n3161) );
  INVX2 U2237 ( .A(n2331), .Y(n2332) );
  OR2X2 U2238 ( .A(n3662), .B(n2332), .Y(n3163) );
  INVX2 U2239 ( .A(n2316), .Y(n2317) );
  INVX4 U2240 ( .A(n2481), .Y(n2482) );
  OR2X2 U2241 ( .A(\sub_x_1100_2/A[6] ), .B(\lt_x_1100_4/B[6] ), .Y(n2446) );
  INVX4 U2242 ( .A(n2479), .Y(n2480) );
  OR2X2 U2243 ( .A(\sub_x_1100_2/A[7] ), .B(\sub_x_1100_2/n227 ), .Y(n2336) );
  INVX2 U2244 ( .A(n3527), .Y(n3526) );
  OR2X2 U2245 ( .A(\sub_x_1100_2/B[4] ), .B(aluOperand1[4]), .Y(n3177) );
  INVX2 U2246 ( .A(n3177), .Y(n3178) );
  INVX2 U2247 ( .A(n3666), .Y(n3667) );
  INVX2 U2248 ( .A(n3198), .Y(n3199) );
  OR2X2 U2249 ( .A(n2060), .B(\lt_x_1100_4/B[15] ), .Y(n2313) );
  INVX2 U2250 ( .A(n3519), .Y(n3518) );
  INVX4 U2251 ( .A(n3202), .Y(n3203) );
  INVX2 U2252 ( .A(n3204), .Y(n3205) );
  INVX2 U2253 ( .A(n2322), .Y(n2323) );
  INVX4 U2254 ( .A(n3528), .Y(n3529) );
  INVX2 U2255 ( .A(n3289), .Y(n3288) );
  OR2X2 U2256 ( .A(aluOperation[3]), .B(aluOperation[0]), .Y(n3166) );
  INVX4 U2257 ( .A(n2337), .Y(n2338) );
  BUFX4 U2258 ( .A(aluResult[30]), .Y(n2225) );
  INVX2 U2259 ( .A(n1818), .Y(n3906) );
  INVX1 U2260 ( .A(n2691), .Y(n2227) );
  INVX1 U2261 ( .A(n2841), .Y(n2235) );
  BUFX4 U2262 ( .A(\ashr_1100_6/SH[0] ), .Y(n4022) );
  BUFX2 U2263 ( .A(n3795), .Y(n3382) );
  BUFX2 U2264 ( .A(n3796), .Y(n3381) );
  BUFX2 U2265 ( .A(n3935), .Y(n3476) );
  BUFX2 U2266 ( .A(n3934), .Y(n3472) );
  BUFX2 U2267 ( .A(n3938), .Y(n3477) );
  INVX1 U2268 ( .A(n2689), .Y(n2228) );
  INVX1 U2269 ( .A(n3235), .Y(n2229) );
  INVX8 U2270 ( .A(n4022), .Y(n2230) );
  INVX1 U2271 ( .A(n2925), .Y(n2231) );
  INVX1 U2272 ( .A(n2496), .Y(n2232) );
  INVX1 U2273 ( .A(\lt_x_1100_4/B[10] ), .Y(n2233) );
  INVX1 U2274 ( .A(n2688), .Y(n2234) );
  INVX8 U2275 ( .A(n2239), .Y(n2236) );
  INVX2 U2276 ( .A(n3709), .Y(n2240) );
  INVX2 U2277 ( .A(n3704), .Y(n2241) );
  BUFX2 U2278 ( .A(n941), .Y(n3085) );
  BUFX2 U2279 ( .A(n4199), .Y(n2492) );
  BUFX2 U2280 ( .A(n4204), .Y(n2493) );
  AND2X1 U2281 ( .A(n2756), .B(n2239), .Y(n2307) );
  AND2X1 U2282 ( .A(n2748), .B(n2239), .Y(n2339) );
  AND2X1 U2283 ( .A(n2760), .B(n2239), .Y(n2348) );
  BUFX2 U2284 ( .A(n3776), .Y(n2246) );
  BUFX2 U2285 ( .A(n3737), .Y(n2248) );
  BUFX2 U2286 ( .A(n3742), .Y(n2247) );
  BUFX2 U2287 ( .A(n3744), .Y(n2244) );
  BUFX2 U2288 ( .A(n3743), .Y(n2245) );
  AND2X1 U2289 ( .A(\sub_x_1100_2/A[0] ), .B(n2230), .Y(n2899) );
  AND2X1 U2290 ( .A(\sub_x_1100_2/A[31] ), .B(n3685), .Y(n2905) );
  BUFX2 U2291 ( .A(n3773), .Y(n2249) );
  BUFX2 U2292 ( .A(n3775), .Y(n2255) );
  INVX1 U2293 ( .A(n2277), .Y(n2237) );
  AND2X1 U2294 ( .A(n1138), .B(n1140), .Y(n3502) );
  AND2X1 U2295 ( .A(n4334), .B(n4333), .Y(n2503) );
  AND2X1 U2296 ( .A(n1138), .B(n1141), .Y(n3508) );
  BUFX2 U2297 ( .A(n933), .Y(n3082) );
  BUFX2 U2298 ( .A(n913), .Y(n3078) );
  BUFX2 U2299 ( .A(n917), .Y(n3080) );
  BUFX2 U2300 ( .A(n4187), .Y(n2802) );
  BUFX2 U2301 ( .A(n3947), .Y(n2980) );
  BUFX2 U2302 ( .A(n3869), .Y(n3326) );
  BUFX2 U2303 ( .A(n3899), .Y(n3330) );
  BUFX2 U2304 ( .A(n3844), .Y(n3405) );
  BUFX2 U2305 ( .A(n3855), .Y(n3411) );
  BUFX2 U2306 ( .A(n3835), .Y(n3271) );
  BUFX2 U2307 ( .A(n4192), .Y(n2831) );
  BUFX2 U2308 ( .A(n4186), .Y(n2830) );
  BUFX2 U2309 ( .A(\sub_x_1100_2/n94 ), .Y(n2686) );
  BUFX2 U2310 ( .A(\add_x_1100_1/n75 ), .Y(n2681) );
  BUFX2 U2311 ( .A(n4202), .Y(n2635) );
  INVX1 U2312 ( .A(n2899), .Y(n2900) );
  INVX1 U2313 ( .A(n2905), .Y(n2906) );
  AND2X1 U2314 ( .A(n3211), .B(\add_x_1100_1/n195 ), .Y(n3109) );
  BUFX2 U2315 ( .A(n4197), .Y(n2633) );
  AND2X1 U2316 ( .A(n2253), .B(n3238), .Y(n2819) );
  INVX1 U2317 ( .A(n3522), .Y(n3523) );
  INVX1 U2318 ( .A(n3544), .Y(n3545) );
  BUFX2 U2319 ( .A(n3769), .Y(n2917) );
  BUFX2 U2320 ( .A(n4184), .Y(n2961) );
  BUFX2 U2321 ( .A(n3785), .Y(n3238) );
  BUFX2 U2322 ( .A(n4190), .Y(n2962) );
  INVX8 U2323 ( .A(n3906), .Y(n2238) );
  BUFX2 U2324 ( .A(n2286), .Y(n3909) );
  INVX1 U2325 ( .A(n3179), .Y(n3180) );
  AND2X1 U2326 ( .A(aluOperand1[21]), .B(n3245), .Y(n2497) );
  AND2X1 U2327 ( .A(aluOperand1[25]), .B(n3241), .Y(n2993) );
  AND2X1 U2328 ( .A(aluOperand1[19]), .B(n3247), .Y(n2690) );
  INVX1 U2329 ( .A(\lt_x_1100_4/B[17] ), .Y(n2257) );
  INVX1 U2330 ( .A(\lt_x_1100_4/B[16] ), .Y(n2263) );
  INVX8 U2331 ( .A(n3907), .Y(n2239) );
  INVX1 U2332 ( .A(n2283), .Y(n2242) );
  AND2X2 U2333 ( .A(n3720), .B(n4324), .Y(n2490) );
  INVX1 U2334 ( .A(n3302), .Y(n3303) );
  INVX1 U2335 ( .A(n3186), .Y(n3187) );
  INVX1 U2336 ( .A(n3505), .Y(n3506) );
  BUFX2 U2337 ( .A(n965), .Y(n3093) );
  BUFX2 U2338 ( .A(n961), .Y(n3092) );
  BUFX2 U2339 ( .A(n4282), .Y(n2813) );
  BUFX2 U2340 ( .A(n957), .Y(n3090) );
  BUFX2 U2341 ( .A(n959), .Y(n3091) );
  BUFX2 U2342 ( .A(n4275), .Y(n2812) );
  BUFX2 U2343 ( .A(n4267), .Y(n2811) );
  BUFX2 U2344 ( .A(n4252), .Y(n2809) );
  BUFX2 U2345 ( .A(n953), .Y(n3089) );
  BUFX2 U2346 ( .A(n4260), .Y(n2810) );
  BUFX2 U2347 ( .A(n945), .Y(n3086) );
  OR2X1 U2348 ( .A(n2805), .B(n2311), .Y(n2310) );
  BUFX2 U2349 ( .A(n4245), .Y(n2808) );
  BUFX2 U2350 ( .A(n4237), .Y(n2807) );
  BUFX2 U2351 ( .A(n4227), .Y(n2806) );
  OR2X1 U2352 ( .A(n3020), .B(n2939), .Y(n2311) );
  BUFX2 U2353 ( .A(n4211), .Y(n2804) );
  AND2X1 U2354 ( .A(n2492), .B(n2634), .Y(n921) );
  AND2X1 U2355 ( .A(n2493), .B(n2798), .Y(n923) );
  BUFX2 U2356 ( .A(n4244), .Y(n2834) );
  BUFX2 U2357 ( .A(n4236), .Y(n2833) );
  BUFX2 U2358 ( .A(n4193), .Y(n2803) );
  BUFX2 U2359 ( .A(n4251), .Y(n2835) );
  AND2X1 U2360 ( .A(aluOperation[3]), .B(n2632), .Y(n2939) );
  BUFX2 U2361 ( .A(n4281), .Y(n2839) );
  BUFX2 U2362 ( .A(\sub_x_1100_2/n84 ), .Y(n3062) );
  BUFX2 U2363 ( .A(n4266), .Y(n2837) );
  BUFX2 U2364 ( .A(n4198), .Y(n2634) );
  BUFX2 U2365 ( .A(\arithmetic_logic_unit/N298 ), .Y(n2632) );
  BUFX2 U2366 ( .A(n4274), .Y(n2838) );
  BUFX2 U2367 ( .A(n4226), .Y(n2832) );
  BUFX2 U2368 ( .A(\add_x_1100_1/n80 ), .Y(n3058) );
  INVX1 U2369 ( .A(n2368), .Y(n2369) );
  BUFX2 U2370 ( .A(n4259), .Y(n2836) );
  BUFX2 U2371 ( .A(\sub_x_1100_2/n99 ), .Y(n3063) );
  BUFX2 U2372 ( .A(\add_x_1100_1/n95 ), .Y(n3059) );
  BUFX2 U2373 ( .A(n4288), .Y(n2840) );
  AND2X1 U2374 ( .A(n4293), .B(n2745), .Y(n2368) );
  OR2X1 U2375 ( .A(n3907), .B(n3327), .Y(n2391) );
  BUFX2 U2376 ( .A(n3898), .Y(n3329) );
  AND2X1 U2377 ( .A(n2373), .B(n4293), .Y(n3017) );
  BUFX2 U2378 ( .A(n3998), .Y(n3333) );
  BUFX2 U2379 ( .A(n3875), .Y(n3327) );
  BUFX2 U2380 ( .A(n3962), .Y(n2984) );
  AND2X1 U2381 ( .A(n2498), .B(n2633), .Y(n2823) );
  BUFX2 U2382 ( .A(n4003), .Y(n2760) );
  BUFX2 U2383 ( .A(n4004), .Y(n3334) );
  BUFX2 U2384 ( .A(n3997), .Y(n2759) );
  BUFX2 U2385 ( .A(n3894), .Y(n3358) );
  BUFX2 U2386 ( .A(n3845), .Y(n2750) );
  BUFX2 U2387 ( .A(n3881), .Y(n2756) );
  BUFX2 U2388 ( .A(n3963), .Y(n3361) );
  BUFX2 U2389 ( .A(n3874), .Y(n2755) );
  AND2X1 U2390 ( .A(n2500), .B(n2635), .Y(n2825) );
  BUFX2 U2391 ( .A(n3868), .Y(n2754) );
  BUFX2 U2392 ( .A(n3856), .Y(n2752) );
  OR2X1 U2393 ( .A(n2236), .B(n3350), .Y(n2867) );
  BUFX2 U2394 ( .A(n3987), .Y(n2758) );
  BUFX2 U2395 ( .A(n3850), .Y(n2751) );
  BUFX2 U2396 ( .A(n3863), .Y(n2753) );
  BUFX2 U2397 ( .A(n3979), .Y(n3331) );
  BUFX2 U2398 ( .A(n4008), .Y(n3335) );
  OR2X1 U2399 ( .A(n3907), .B(n3344), .Y(n2344) );
  BUFX2 U2400 ( .A(n3992), .Y(n3362) );
  AND2X1 U2401 ( .A(n3908), .B(n3299), .Y(n3346) );
  BUFX2 U2402 ( .A(n3823), .Y(n2748) );
  BUFX2 U2403 ( .A(n3886), .Y(n3356) );
  BUFX2 U2404 ( .A(n3948), .Y(n3359) );
  BUFX2 U2405 ( .A(\sub_x_1100_2/n124 ), .Y(n3064) );
  OR2X1 U2406 ( .A(n3907), .B(n3340), .Y(n2372) );
  BUFX2 U2407 ( .A(n3840), .Y(n2749) );
  BUFX2 U2408 ( .A(n3890), .Y(n3357) );
  BUFX2 U2409 ( .A(n3925), .Y(n2757) );
  BUFX2 U2410 ( .A(n3832), .Y(n3299) );
  BUFX2 U2411 ( .A(\sub_x_1100_2/n155 ), .Y(n3065) );
  BUFX2 U2412 ( .A(\sub_x_1100_2/n150 ), .Y(n3516) );
  BUFX2 U2413 ( .A(n4007), .Y(n3281) );
  BUFX2 U2414 ( .A(n3879), .Y(n2979) );
  BUFX2 U2415 ( .A(n3873), .Y(n3420) );
  BUFX2 U2416 ( .A(n4012), .Y(n3495) );
  BUFX2 U2417 ( .A(n4013), .Y(n3492) );
  BUFX2 U2418 ( .A(n3867), .Y(n3417) );
  BUFX2 U2419 ( .A(n3885), .Y(n3426) );
  BUFX2 U2420 ( .A(n3872), .Y(n2977) );
  BUFX2 U2421 ( .A(n4001), .Y(n2988) );
  BUFX2 U2422 ( .A(n3827), .Y(n3268) );
  BUFX2 U2423 ( .A(n3851), .Y(n3272) );
  BUFX2 U2424 ( .A(n3849), .Y(n3408) );
  BUFX2 U2425 ( .A(n3995), .Y(n2987) );
  BUFX2 U2426 ( .A(n3986), .Y(n3482) );
  BUFX2 U2427 ( .A(n3866), .Y(n2976) );
  BUFX2 U2428 ( .A(n3972), .Y(n3375) );
  BUFX2 U2429 ( .A(n3831), .Y(n3269) );
  BUFX2 U2430 ( .A(n3970), .Y(n3491) );
  BUFX2 U2431 ( .A(n4009), .Y(n3460) );
  BUFX2 U2432 ( .A(n3841), .Y(n3371) );
  BUFX2 U2433 ( .A(n3961), .Y(n2983) );
  BUFX2 U2434 ( .A(n3991), .Y(n3484) );
  BUFX2 U2435 ( .A(n4002), .Y(n3280) );
  BUFX2 U2436 ( .A(n3839), .Y(n3402) );
  AND2X1 U2437 ( .A(n3908), .B(n3301), .Y(n3351) );
  BUFX2 U2438 ( .A(n3978), .Y(n3468) );
  BUFX2 U2439 ( .A(n3969), .Y(n3490) );
  BUFX2 U2440 ( .A(n3893), .Y(n3432) );
  BUFX2 U2441 ( .A(n3985), .Y(n2986) );
  BUFX2 U2442 ( .A(n3836), .Y(n3370) );
  BUFX2 U2443 ( .A(n3854), .Y(n2974) );
  BUFX2 U2444 ( .A(n3862), .Y(n3414) );
  BUFX2 U2445 ( .A(n3861), .Y(n2975) );
  BUFX2 U2446 ( .A(n3889), .Y(n3429) );
  BUFX2 U2447 ( .A(n3953), .Y(n3275) );
  BUFX2 U2448 ( .A(n3857), .Y(n3273) );
  AND2X1 U2449 ( .A(n3908), .B(n3300), .Y(n3349) );
  BUFX2 U2450 ( .A(n3966), .Y(n3483) );
  BUFX2 U2451 ( .A(n3973), .Y(n3336) );
  BUFX2 U2452 ( .A(n4010), .Y(n3453) );
  BUFX2 U2453 ( .A(n3846), .Y(n3372) );
  BUFX2 U2454 ( .A(n3971), .Y(n3374) );
  AND2X1 U2455 ( .A(n3292), .B(n3908), .Y(n3367) );
  BUFX2 U2456 ( .A(n3956), .Y(n3301) );
  BUFX2 U2457 ( .A(\add_x_1100_1/n120 ), .Y(n3060) );
  BUFX2 U2458 ( .A(n3954), .Y(n3300) );
  AND2X1 U2459 ( .A(n3294), .B(n3908), .Y(n3369) );
  BUFX2 U2460 ( .A(\add_x_1100_1/n151 ), .Y(n3061) );
  BUFX2 U2461 ( .A(\add_x_1100_1/n146 ), .Y(n3513) );
  AND2X1 U2462 ( .A(n3290), .B(n3908), .Y(n3339) );
  BUFX2 U2463 ( .A(n3951), .Y(n3487) );
  BUFX2 U2464 ( .A(n3945), .Y(n3478) );
  BUFX2 U2465 ( .A(n3814), .Y(n3394) );
  BUFX2 U2466 ( .A(n3928), .Y(n3456) );
  BUFX2 U2467 ( .A(n3779), .Y(n2892) );
  BUFX2 U2468 ( .A(n3984), .Y(n2985) );
  BUFX2 U2469 ( .A(n3811), .Y(n3391) );
  BUFX2 U2470 ( .A(n3812), .Y(n3355) );
  BUFX2 U2471 ( .A(n3958), .Y(n3488) );
  BUFX2 U2472 ( .A(n3946), .Y(n3475) );
  BUFX2 U2473 ( .A(n3793), .Y(n3380) );
  BUFX2 U2474 ( .A(n3994), .Y(n3494) );
  BUFX2 U2475 ( .A(n4005), .Y(n3500) );
  BUFX2 U2476 ( .A(n3990), .Y(n3459) );
  BUFX2 U2477 ( .A(n4006), .Y(n3481) );
  BUFX2 U2478 ( .A(n3741), .Y(n3239) );
  BUFX2 U2479 ( .A(n3747), .Y(n3379) );
  BUFX2 U2480 ( .A(n3834), .Y(n3410) );
  BUFX2 U2481 ( .A(n3826), .Y(n3404) );
  BUFX2 U2482 ( .A(n3941), .Y(n3466) );
  BUFX2 U2483 ( .A(n3871), .Y(n3431) );
  BUFX2 U2484 ( .A(n3810), .Y(n3387) );
  BUFX2 U2485 ( .A(n3818), .Y(n3397) );
  BUFX2 U2486 ( .A(n4000), .Y(n3467) );
  BUFX2 U2487 ( .A(n3950), .Y(n3360) );
  BUFX2 U2488 ( .A(n3993), .Y(n3498) );
  BUFX2 U2489 ( .A(n3853), .Y(n3422) );
  BUFX2 U2490 ( .A(n3815), .Y(n3395) );
  BUFX2 U2491 ( .A(n3820), .Y(n3398) );
  BUFX2 U2492 ( .A(n3843), .Y(n3416) );
  BUFX2 U2493 ( .A(n3960), .Y(n2982) );
  BUFX2 U2494 ( .A(n3807), .Y(n3384) );
  BUFX2 U2495 ( .A(n3830), .Y(n3407) );
  BUFX2 U2496 ( .A(n3892), .Y(n3440) );
  BUFX2 U2497 ( .A(n3819), .Y(n3399) );
  BUFX2 U2498 ( .A(n3865), .Y(n3428) );
  BUFX2 U2499 ( .A(n3952), .Y(n3486) );
  BUFX2 U2500 ( .A(n3888), .Y(n3438) );
  BUFX2 U2501 ( .A(n3878), .Y(n3434) );
  BUFX2 U2502 ( .A(n3848), .Y(n3419) );
  BUFX2 U2503 ( .A(n3949), .Y(n3485) );
  BUFX2 U2504 ( .A(n3808), .Y(n3354) );
  BUFX2 U2505 ( .A(n3822), .Y(n3401) );
  BUFX2 U2506 ( .A(n3838), .Y(n3413) );
  BUFX2 U2507 ( .A(n3860), .Y(n3425) );
  BUFX2 U2508 ( .A(n3816), .Y(n3270) );
  BUFX2 U2509 ( .A(n3877), .Y(n2978) );
  BUFX2 U2510 ( .A(n3884), .Y(n3436) );
  BUFX2 U2511 ( .A(n3989), .Y(n3463) );
  BUFX2 U2512 ( .A(n3999), .Y(n3499) );
  BUFX2 U2513 ( .A(n3965), .Y(n3550) );
  BUFX2 U2514 ( .A(n3944), .Y(n3276) );
  BUFX2 U2515 ( .A(n3782), .Y(n3325) );
  BUFX2 U2516 ( .A(n3926), .Y(n3449) );
  BUFX2 U2517 ( .A(n3730), .Y(n2829) );
  BUFX2 U2518 ( .A(n3942), .Y(n3465) );
  BUFX2 U2519 ( .A(n3929), .Y(n3452) );
  BUFX2 U2520 ( .A(n3940), .Y(n3274) );
  BUFX2 U2521 ( .A(n3927), .Y(n3446) );
  BUFX2 U2522 ( .A(n4208), .Y(n2963) );
  BUFX2 U2523 ( .A(n3930), .Y(n3469) );
  BUFX2 U2524 ( .A(n3933), .Y(n3473) );
  BUFX2 U2525 ( .A(n3802), .Y(n3389) );
  BUFX2 U2526 ( .A(n3870), .Y(n3435) );
  BUFX2 U2527 ( .A(n3859), .Y(n3430) );
  BUFX2 U2528 ( .A(n3891), .Y(n3442) );
  BUFX2 U2529 ( .A(n3883), .Y(n3439) );
  BUFX2 U2530 ( .A(n3976), .Y(n3464) );
  BUFX2 U2531 ( .A(n3798), .Y(n3385) );
  BUFX2 U2532 ( .A(n3847), .Y(n3424) );
  BUFX2 U2533 ( .A(n3837), .Y(n3418) );
  BUFX2 U2534 ( .A(n3801), .Y(n3363) );
  BUFX2 U2535 ( .A(n3829), .Y(n3412) );
  BUFX2 U2536 ( .A(n3821), .Y(n3406) );
  BUFX2 U2537 ( .A(n3813), .Y(n3400) );
  BUFX2 U2538 ( .A(n3803), .Y(n3388) );
  BUFX2 U2539 ( .A(n3806), .Y(n3393) );
  BUFX2 U2540 ( .A(n3977), .Y(n3462) );
  BUFX2 U2541 ( .A(n3804), .Y(n3392) );
  BUFX2 U2542 ( .A(n3959), .Y(n2981) );
  BUFX2 U2543 ( .A(n3805), .Y(n3390) );
  BUFX2 U2544 ( .A(n3980), .Y(n3496) );
  BUFX2 U2545 ( .A(n3974), .Y(n3461) );
  BUFX2 U2546 ( .A(n3833), .Y(n3415) );
  BUFX2 U2547 ( .A(n3876), .Y(n3437) );
  BUFX2 U2548 ( .A(n3887), .Y(n3441) );
  AND2X1 U2549 ( .A(n2255), .B(n3168), .Y(n3312) );
  BUFX2 U2550 ( .A(n3800), .Y(n3386) );
  BUFX2 U2551 ( .A(n3817), .Y(n3403) );
  BUFX2 U2552 ( .A(n3852), .Y(n3427) );
  BUFX2 U2553 ( .A(n3864), .Y(n3433) );
  BUFX2 U2554 ( .A(n3957), .Y(n3480) );
  BUFX2 U2555 ( .A(n3923), .Y(n3455) );
  BUFX2 U2556 ( .A(n3937), .Y(n3479) );
  BUFX2 U2557 ( .A(n3825), .Y(n3409) );
  BUFX2 U2558 ( .A(n3809), .Y(n3396) );
  BUFX2 U2559 ( .A(n3922), .Y(n3457) );
  BUFX2 U2560 ( .A(n3920), .Y(n3454) );
  BUFX2 U2561 ( .A(n3975), .Y(n3458) );
  BUFX2 U2562 ( .A(n3981), .Y(n3493) );
  BUFX2 U2563 ( .A(n3799), .Y(n3383) );
  BUFX2 U2564 ( .A(n3983), .Y(n3497) );
  BUFX2 U2565 ( .A(n3797), .Y(n3364) );
  BUFX2 U2566 ( .A(n3943), .Y(n3365) );
  BUFX2 U2567 ( .A(n3917), .Y(n3445) );
  BUFX2 U2568 ( .A(n3913), .Y(n3444) );
  BUFX2 U2569 ( .A(n3916), .Y(n3447) );
  BUFX2 U2570 ( .A(n3914), .Y(n3443) );
  BUFX2 U2571 ( .A(n3912), .Y(n3373) );
  BUFX2 U2572 ( .A(n3919), .Y(n3448) );
  BUFX2 U2573 ( .A(n3918), .Y(n3450) );
  BUFX2 U2574 ( .A(n3921), .Y(n3451) );
  AND2X1 U2575 ( .A(n2232), .B(n3170), .Y(n2821) );
  BUFX2 U2576 ( .A(\sub_x_1100_2/n79 ), .Y(n2685) );
  AND2X1 U2577 ( .A(n2232), .B(n3169), .Y(n2817) );
  BUFX2 U2578 ( .A(n3770), .Y(n2889) );
  AND2X1 U2579 ( .A(n3157), .B(n3678), .Y(n3637) );
  AND2X1 U2580 ( .A(n2161), .B(n3681), .Y(n3633) );
  AND2X1 U2581 ( .A(n2143), .B(n3679), .Y(n3635) );
  BUFX2 U2582 ( .A(n3729), .Y(n2746) );
  BUFX2 U2583 ( .A(n3774), .Y(n2989) );
  BUFX2 U2584 ( .A(n3784), .Y(n2744) );
  BUFX2 U2585 ( .A(n3788), .Y(n2898) );
  BUFX2 U2586 ( .A(n3783), .Y(n2896) );
  BUFX2 U2587 ( .A(n3789), .Y(n2894) );
  BUFX2 U2588 ( .A(n3745), .Y(n3169) );
  BUFX2 U2589 ( .A(n3792), .Y(n3170) );
  BUFX2 U2590 ( .A(n3786), .Y(n2893) );
  BUFX2 U2591 ( .A(n3731), .Y(n3168) );
  INVX1 U2592 ( .A(n2330), .Y(n2250) );
  BUFX2 U2593 ( .A(n1345), .Y(n2765) );
  BUFX2 U2594 ( .A(n1301), .Y(n2787) );
  BUFX2 U2595 ( .A(n1337), .Y(n2769) );
  BUFX2 U2596 ( .A(n1343), .Y(n2766) );
  BUFX2 U2597 ( .A(n4278), .Y(n2972) );
  BUFX2 U2598 ( .A(n1333), .Y(n2771) );
  BUFX2 U2599 ( .A(n1303), .Y(n2786) );
  BUFX2 U2600 ( .A(n1353), .Y(n2761) );
  BUFX2 U2601 ( .A(n1335), .Y(n2770) );
  BUFX2 U2602 ( .A(n1341), .Y(n2767) );
  BUFX2 U2603 ( .A(n1315), .Y(n2780) );
  BUFX2 U2604 ( .A(n4285), .Y(n2973) );
  BUFX2 U2605 ( .A(n1339), .Y(n2768) );
  BUFX2 U2606 ( .A(n1305), .Y(n2785) );
  BUFX2 U2607 ( .A(n1323), .Y(n2776) );
  BUFX2 U2608 ( .A(n1293), .Y(n2791) );
  BUFX2 U2609 ( .A(n1311), .Y(n2782) );
  BUFX2 U2610 ( .A(n1321), .Y(n2777) );
  BUFX2 U2611 ( .A(n1349), .Y(n2763) );
  BUFX2 U2612 ( .A(n1307), .Y(n2784) );
  BUFX2 U2613 ( .A(n1347), .Y(n2764) );
  BUFX2 U2614 ( .A(n1288), .Y(n2792) );
  BUFX2 U2615 ( .A(n1317), .Y(n2779) );
  BUFX2 U2616 ( .A(n1309), .Y(n2783) );
  BUFX2 U2617 ( .A(n1351), .Y(n2762) );
  BUFX2 U2618 ( .A(n1313), .Y(n2781) );
  BUFX2 U2619 ( .A(n1319), .Y(n2778) );
  BUFX2 U2620 ( .A(n1329), .Y(n2773) );
  BUFX2 U2621 ( .A(n1327), .Y(n2774) );
  BUFX2 U2622 ( .A(n1297), .Y(n2789) );
  BUFX2 U2623 ( .A(n1295), .Y(n2790) );
  BUFX2 U2624 ( .A(n1299), .Y(n2788) );
  BUFX2 U2625 ( .A(n1325), .Y(n2775) );
  BUFX2 U2626 ( .A(n1331), .Y(n2772) );
  BUFX2 U2627 ( .A(n3791), .Y(n2895) );
  BUFX2 U2628 ( .A(n3780), .Y(n2743) );
  BUFX2 U2629 ( .A(n4264), .Y(n2970) );
  INVX8 U2630 ( .A(n2238), .Y(n2251) );
  BUFX2 U2631 ( .A(n4233), .Y(n2966) );
  INVX1 U2632 ( .A(n2327), .Y(n2328) );
  BUFX2 U2633 ( .A(n4272), .Y(n2971) );
  INVX1 U2634 ( .A(n2993), .Y(n2252) );
  BUFX2 U2635 ( .A(n3768), .Y(n2916) );
  BUFX2 U2636 ( .A(n4241), .Y(n2967) );
  BUFX2 U2637 ( .A(n4249), .Y(n2968) );
  INVX1 U2638 ( .A(n2497), .Y(n2253) );
  BUFX2 U2639 ( .A(n1310), .Y(n2733) );
  BUFX2 U2640 ( .A(n1324), .Y(n2726) );
  BUFX2 U2641 ( .A(n1294), .Y(n2741) );
  BUFX2 U2642 ( .A(n1352), .Y(n2712) );
  BUFX2 U2643 ( .A(n1316), .Y(n2730) );
  BUFX2 U2644 ( .A(n1314), .Y(n2731) );
  BUFX2 U2645 ( .A(n1308), .Y(n2734) );
  BUFX2 U2646 ( .A(n1306), .Y(n2735) );
  BUFX2 U2647 ( .A(n1350), .Y(n2713) );
  BUFX2 U2648 ( .A(n1322), .Y(n2727) );
  BUFX2 U2649 ( .A(n1289), .Y(n2742) );
  BUFX2 U2650 ( .A(n1348), .Y(n2714) );
  BUFX2 U2651 ( .A(n1320), .Y(n2728) );
  BUFX2 U2652 ( .A(n1318), .Y(n2729) );
  BUFX2 U2653 ( .A(n1332), .Y(n2722) );
  BUFX2 U2654 ( .A(n1298), .Y(n2739) );
  BUFX2 U2655 ( .A(n1300), .Y(n2738) );
  BUFX2 U2656 ( .A(n1334), .Y(n2721) );
  BUFX2 U2657 ( .A(n1340), .Y(n2718) );
  BUFX2 U2658 ( .A(n1342), .Y(n2717) );
  BUFX2 U2659 ( .A(n1302), .Y(n2737) );
  BUFX2 U2660 ( .A(n1344), .Y(n2716) );
  BUFX2 U2661 ( .A(n1336), .Y(n2720) );
  BUFX2 U2662 ( .A(n1346), .Y(n2715) );
  BUFX2 U2663 ( .A(n1338), .Y(n2719) );
  BUFX2 U2664 ( .A(n1326), .Y(n2725) );
  BUFX2 U2665 ( .A(n1312), .Y(n2732) );
  BUFX2 U2666 ( .A(n1328), .Y(n2724) );
  BUFX2 U2667 ( .A(n1296), .Y(n2740) );
  BUFX2 U2668 ( .A(n1354), .Y(n2711) );
  BUFX2 U2669 ( .A(n1330), .Y(n2723) );
  BUFX2 U2670 ( .A(n1304), .Y(n2736) );
  INVX1 U2671 ( .A(n2422), .Y(n2423) );
  AND2X1 U2672 ( .A(n3684), .B(n3683), .Y(n2393) );
  BUFX2 U2673 ( .A(n4224), .Y(n2965) );
  INVX1 U2674 ( .A(n2690), .Y(n2254) );
  BUFX2 U2675 ( .A(n4218), .Y(n2964) );
  BUFX2 U2676 ( .A(n3778), .Y(n2891) );
  BUFX2 U2677 ( .A(n3777), .Y(n2890) );
  INVX1 U2678 ( .A(\sub_x_1100_2/n227 ), .Y(n2293) );
  INVX1 U2679 ( .A(n3712), .Y(\ashr_1100_6/SH[3] ) );
  INVX1 U2680 ( .A(n3665), .Y(n2256) );
  OR2X1 U2681 ( .A(aluOperand1[19]), .B(\lt_x_1100_4/B[19] ), .Y(n2422) );
  INVX1 U2682 ( .A(n3661), .Y(n3662) );
  INVX1 U2683 ( .A(n3705), .Y(n2258) );
  INVX1 U2684 ( .A(\lt_x_1100_4/B[8] ), .Y(n2259) );
  BUFX2 U2685 ( .A(n4261), .Y(n3241) );
  BUFX2 U2686 ( .A(n4253), .Y(n3242) );
  BUFX2 U2687 ( .A(n4246), .Y(n3243) );
  BUFX2 U2688 ( .A(n4291), .Y(n3283) );
  BUFX2 U2689 ( .A(n4238), .Y(n3244) );
  BUFX2 U2690 ( .A(n4229), .Y(n3246) );
  BUFX2 U2691 ( .A(n4286), .Y(n3257) );
  BUFX2 U2692 ( .A(n4230), .Y(n3245) );
  BUFX2 U2693 ( .A(n4279), .Y(n3258) );
  BUFX2 U2694 ( .A(n4268), .Y(n3240) );
  OR2X1 U2695 ( .A(n4329), .B(n4034), .Y(n3713) );
  OR2X1 U2696 ( .A(n2279), .B(n4034), .Y(n3714) );
  BUFX2 U2697 ( .A(n4221), .Y(n3248) );
  BUFX2 U2698 ( .A(n4228), .Y(n3247) );
  BUFX2 U2699 ( .A(n4292), .Y(n3282) );
  OR2X1 U2700 ( .A(n2432), .B(n245), .Y(n3710) );
  BUFX2 U2701 ( .A(n4033), .Y(n2828) );
  OR2X1 U2702 ( .A(n2795), .B(instructionType[2]), .Y(n847) );
  BUFX2 U2703 ( .A(n4045), .Y(n2656) );
  BUFX2 U2704 ( .A(n4047), .Y(n2657) );
  BUFX2 U2705 ( .A(n4039), .Y(n2653) );
  BUFX2 U2706 ( .A(n4037), .Y(n2652) );
  BUFX2 U2707 ( .A(n4043), .Y(n2655) );
  BUFX2 U2708 ( .A(n4041), .Y(n2654) );
  BUFX2 U2709 ( .A(n4049), .Y(n2658) );
  BUFX2 U2710 ( .A(n4051), .Y(n2659) );
  BUFX2 U2711 ( .A(n4053), .Y(n2660) );
  BUFX2 U2712 ( .A(n848), .Y(n4032) );
  BUFX2 U2713 ( .A(n4169), .Y(n2795) );
  BUFX2 U2714 ( .A(n4057), .Y(n2662) );
  INVX1 U2715 ( .A(n2283), .Y(n2265) );
  BUFX2 U2716 ( .A(n555), .Y(n3073) );
  BUFX2 U2717 ( .A(n557), .Y(n3074) );
  AND2X1 U2718 ( .A(aluResultRegister[29]), .B(n4024), .Y(n2999) );
  AND2X1 U2719 ( .A(pc[28]), .B(n2299), .Y(n2934) );
  AND2X1 U2720 ( .A(pc[29]), .B(n2299), .Y(n2932) );
  AND2X1 U2721 ( .A(aluResultRegister[28]), .B(n4024), .Y(n3001) );
  AND2X1 U2722 ( .A(aluResultRegister[30]), .B(n4024), .Y(n2997) );
  AND2X1 U2723 ( .A(pc[30]), .B(n2299), .Y(n2930) );
  AND2X1 U2724 ( .A(aluResultRegister[27]), .B(n4024), .Y(n3003) );
  AND2X1 U2725 ( .A(pc[27]), .B(n2298), .Y(n3631) );
  AND2X1 U2726 ( .A(aluResultRegister[31]), .B(n4024), .Y(n2995) );
  AND2X1 U2727 ( .A(pc[31]), .B(n2299), .Y(n2928) );
  BUFX2 U2728 ( .A(N924), .Y(n3054) );
  BUFX2 U2729 ( .A(n4167), .Y(n2856) );
  BUFX2 U2730 ( .A(n4360), .Y(n3561) );
  BUFX2 U2731 ( .A(n4157), .Y(n2801) );
  AND2X1 U2732 ( .A(n4030), .B(n2295), .Y(n3623) );
  AND2X1 U2733 ( .A(n4030), .B(n2305), .Y(n3617) );
  AND2X1 U2734 ( .A(n4030), .B(n2285), .Y(n3619) );
  AND2X1 U2735 ( .A(n4030), .B(n2294), .Y(n3621) );
  BUFX2 U2736 ( .A(n4156), .Y(n2855) );
  AND2X1 U2737 ( .A(n4030), .B(N1168), .Y(n3599) );
  BUFX2 U2738 ( .A(n551), .Y(n3072) );
  BUFX2 U2739 ( .A(n549), .Y(n3070) );
  AND2X1 U2740 ( .A(n2491), .B(n2799), .Y(n513) );
  AND2X1 U2741 ( .A(n4163), .B(n2638), .Y(n3013) );
  BUFX2 U2742 ( .A(n504), .Y(n3057) );
  AND2X1 U2743 ( .A(n3560), .B(n2648), .Y(n3322) );
  AND2X1 U2744 ( .A(n2502), .B(n2637), .Y(n3155) );
  BUFX2 U2745 ( .A(n4152), .Y(n2992) );
  BUFX2 U2746 ( .A(n4331), .Y(n2793) );
  BUFX2 U2747 ( .A(n1449), .Y(n2638) );
  BUFX2 U2748 ( .A(n4134), .Y(n3296) );
  BUFX2 U2749 ( .A(n4321), .Y(n3045) );
  BUFX2 U2750 ( .A(n4335), .Y(n2637) );
  BUFX2 U2751 ( .A(n4127), .Y(n2491) );
  BUFX2 U2752 ( .A(n4116), .Y(n2796) );
  BUFX2 U2753 ( .A(n4339), .Y(n2857) );
  BUFX2 U2754 ( .A(n4162), .Y(n2960) );
  BUFX2 U2755 ( .A(n4124), .Y(n2879) );
  AND2X1 U2756 ( .A(n2495), .B(n2639), .Y(n3504) );
  BUFX2 U2757 ( .A(n4133), .Y(n3304) );
  BUFX2 U2758 ( .A(n4144), .Y(n3554) );
  BUFX2 U2759 ( .A(n977), .Y(n3376) );
  BUFX2 U2760 ( .A(n4137), .Y(n2800) );
  BUFX2 U2761 ( .A(n1426), .Y(n2923) );
  BUFX2 U2762 ( .A(n982), .Y(n2639) );
  AND2X1 U2763 ( .A(n4328), .B(n2636), .Y(n2827) );
  AND2X1 U2764 ( .A(n1144), .B(n2455), .Y(n4159) );
  BUFX2 U2765 ( .A(n4114), .Y(n2922) );
  INVX1 U2766 ( .A(n2424), .Y(n2267) );
  BUFX2 U2767 ( .A(n4132), .Y(n3039) );
  AND2X1 U2768 ( .A(n2494), .B(n4334), .Y(n2886) );
  AND2X1 U2769 ( .A(n4373), .B(n4168), .Y(n3005) );
  BUFX2 U2770 ( .A(n4327), .Y(n2636) );
  INVX1 U2771 ( .A(n2408), .Y(n2268) );
  BUFX2 U2772 ( .A(n980), .Y(n3517) );
  BUFX2 U2773 ( .A(n981), .Y(n2495) );
  AND2X1 U2774 ( .A(n3559), .B(n2437), .Y(n3049) );
  BUFX2 U2775 ( .A(n4375), .Y(n2494) );
  INVX1 U2776 ( .A(n2486), .Y(n2269) );
  INVX1 U2777 ( .A(n3167), .Y(n2270) );
  BUFX2 U2778 ( .A(n4128), .Y(n2913) );
  BUFX2 U2779 ( .A(n1427), .Y(n3530) );
  BUFX2 U2780 ( .A(n4150), .Y(n3549) );
  AND2X1 U2781 ( .A(n4120), .B(n3674), .Y(n4112) );
  INVX1 U2782 ( .A(n2363), .Y(n2271) );
  INVX1 U2783 ( .A(opcode[6]), .Y(n2272) );
  INVX1 U2784 ( .A(aluZeroRegister), .Y(n2289) );
  AND2X2 U2785 ( .A(\lt_x_1100_4/B[8] ), .B(n2743), .Y(n2689) );
  INVX4 U2786 ( .A(n3706), .Y(\ashr_1100_6/SH[0] ) );
  INVX1 U2787 ( .A(n2325), .Y(n2273) );
  INVX2 U2788 ( .A(n4091), .Y(n4024) );
  BUFX2 U2789 ( .A(aluOperand1[4]), .Y(\sub_x_1100_2/A[4] ) );
  AND2X2 U2790 ( .A(aluOperand1[3]), .B(n3712), .Y(n3235) );
  OR2X2 U2791 ( .A(n3712), .B(aluOperand1[3]), .Y(n3666) );
  OR2X2 U2792 ( .A(n2469), .B(n2260), .Y(n2461) );
  OR2X2 U2793 ( .A(n2462), .B(n2256), .Y(n2451) );
  INVX1 U2794 ( .A(aluSrcA[1]), .Y(n2274) );
  AND2X2 U2795 ( .A(n2261), .B(\sub_x_1100_2/A[5] ), .Y(n3234) );
  AND2X2 U2796 ( .A(\sub_x_1100_2/A[2] ), .B(n3707), .Y(n3544) );
  BUFX2 U2797 ( .A(aluOperand1[0]), .Y(\sub_x_1100_2/A[0] ) );
  OAI21X1 U2798 ( .A(n2421), .B(n3512), .C(n3194), .Y(n2275) );
  INVX2 U2799 ( .A(n3675), .Y(n4366) );
  BUFX2 U2800 ( .A(aluOperand1[10]), .Y(\sub_x_1100_2/A[10] ) );
  AND2X2 U2801 ( .A(\lt_x_1100_4/B[9] ), .B(n2470), .Y(n3204) );
  INVX1 U2802 ( .A(n3313), .Y(n2276) );
  AND2X2 U2803 ( .A(\sub_x_1100_2/n228 ), .B(\sub_x_1100_2/A[6] ), .Y(n3668)
         );
  OR2X2 U2804 ( .A(\sub_x_1100_2/A[6] ), .B(\sub_x_1100_2/n228 ), .Y(n3539) );
  AND2X2 U2805 ( .A(n2292), .B(\sub_x_1100_2/A[6] ), .Y(n2481) );
  OR2X2 U2806 ( .A(aluSrcA[0]), .B(aluSrcA[1]), .Y(n2277) );
  AND2X2 U2807 ( .A(aluSrcA[0]), .B(n1852), .Y(n2278) );
  BUFX2 U2808 ( .A(opcode[2]), .Y(n2279) );
  INVX1 U2809 ( .A(n2283), .Y(n2281) );
  INVX1 U2810 ( .A(n2283), .Y(n2284) );
  OR2X2 U2811 ( .A(aluSrcB[0]), .B(aluSrcB[1]), .Y(n2350) );
  BUFX2 U2812 ( .A(N1198), .Y(n2285) );
  AND2X2 U2813 ( .A(n4168), .B(n4109), .Y(n2379) );
  INVX2 U2814 ( .A(n3535), .Y(n2438) );
  OR2X2 U2815 ( .A(n3670), .B(aluOperand1[4]), .Y(n3179) );
  AND2X2 U2816 ( .A(aluOperand1[4]), .B(n3670), .Y(n3527) );
  AND2X2 U2817 ( .A(pc[0]), .B(n2297), .Y(n3703) );
  AND2X2 U2818 ( .A(n2313), .B(n2314), .Y(n2287) );
  AND2X2 U2819 ( .A(n3724), .B(n3726), .Y(n4322) );
  OR2X2 U2820 ( .A(n2379), .B(n3558), .Y(n2288) );
  MUX2X1 U2821 ( .B(\funct3[0] ), .A(n2271), .S(n2289), .Y(n4139) );
  BUFX2 U2822 ( .A(n3286), .Y(n2291) );
  AND2X2 U2823 ( .A(aluOperand1[0]), .B(\ashr_1100_6/SH[0] ), .Y(n2329) );
  OR2X2 U2824 ( .A(n3706), .B(aluOperand1[0]), .Y(n3655) );
  AND2X1 U2825 ( .A(n2215), .B(RS2[0]), .Y(n2376) );
  AND2X1 U2826 ( .A(n2284), .B(RS2[3]), .Y(n2351) );
  BUFX2 U2827 ( .A(\lt_x_1100_4/B[6] ), .Y(n2292) );
  OR2X2 U2828 ( .A(n3705), .B(aluOperand1[1]), .Y(n3289) );
  AND2X2 U2829 ( .A(aluOperand1[1]), .B(n3705), .Y(n3237) );
  AND2X2 U2830 ( .A(n3250), .B(\sub_x_1100_2/A[14] ), .Y(n3522) );
  AND2X2 U2831 ( .A(n3249), .B(\sub_x_1100_2/A[14] ), .Y(n3519) );
  BUFX2 U2832 ( .A(N1201), .Y(n2294) );
  AND2X2 U2833 ( .A(\lt_x_1100_4/B[10] ), .B(aluOperand1[10]), .Y(n3256) );
  BUFX2 U2834 ( .A(N1204), .Y(n2295) );
  OR2X2 U2835 ( .A(n3707), .B(\sub_x_1100_2/A[2] ), .Y(n3528) );
  AND2X2 U2836 ( .A(RS1[0]), .B(n2278), .Y(n3702) );
  AND2X2 U2837 ( .A(\lt_x_1100_4/B[5] ), .B(aluOperand1[5]), .Y(n3209) );
  INVX1 U2838 ( .A(n2319), .Y(n2296) );
  OR2X2 U2839 ( .A(aluOperand1[7]), .B(\lt_x_1100_4/B[7] ), .Y(n2479) );
  AND2X2 U2840 ( .A(\lt_x_1100_4/B[7] ), .B(aluOperand1[7]), .Y(n3207) );
  INVX8 U2841 ( .A(\ashr_1100_6/SH[1] ), .Y(n3910) );
  OR2X2 U2842 ( .A(\sub_x_1100_2/A[8] ), .B(n2259), .Y(n3665) );
  INVX4 U2843 ( .A(n2468), .Y(n2469) );
  AND2X2 U2844 ( .A(n3251), .B(\sub_x_1100_2/A[12] ), .Y(n3525) );
  BUFX4 U2845 ( .A(aluOperand1[12]), .Y(\sub_x_1100_2/A[12] ) );
  AND2X2 U2846 ( .A(\lt_x_1100_4/B[11] ), .B(aluOperand1[11]), .Y(n3202) );
  INVX1 U2847 ( .A(n2390), .Y(n2297) );
  INVX1 U2848 ( .A(n2277), .Y(n2299) );
  INVX1 U2849 ( .A(n2390), .Y(n2300) );
  INVX1 U2850 ( .A(n2390), .Y(n2301) );
  INVX1 U2851 ( .A(n2277), .Y(n2303) );
  INVX1 U2852 ( .A(n2277), .Y(n2304) );
  OR2X2 U2853 ( .A(aluSrcA[1]), .B(aluSrcA[0]), .Y(n2390) );
  BUFX2 U2854 ( .A(N1195), .Y(n2305) );
  INVX8 U2855 ( .A(n4025), .Y(n2306) );
  BUFX4 U2856 ( .A(aluOperand1[14]), .Y(\sub_x_1100_2/A[14] ) );
  OR2X2 U2857 ( .A(n2270), .B(opcode[5]), .Y(n4330) );
  INVX1 U2858 ( .A(n2307), .Y(n2308) );
  OR2X2 U2859 ( .A(\ashr_1100_6/SH[3] ), .B(aluOperand1[3]), .Y(n2312) );
  OR2X2 U2860 ( .A(\sub_x_1100_2/A[14] ), .B(n3249), .Y(n2314) );
  OR2X2 U2861 ( .A(\sub_x_1100_2/A[12] ), .B(\lt_x_1100_4/B[12] ), .Y(n2315)
         );
  AND2X2 U2862 ( .A(\lt_x_1100_4/B[12] ), .B(\sub_x_1100_2/A[12] ), .Y(n2316)
         );
  AND2X2 U2863 ( .A(n2296), .B(n2410), .Y(n2318) );
  OR2X2 U2864 ( .A(n3532), .B(n2453), .Y(n2319) );
  OR2X2 U2865 ( .A(\lt_x_1100_4/B[11] ), .B(aluOperand1[11]), .Y(n2320) );
  OR2X2 U2866 ( .A(aluOperand1[10]), .B(\lt_x_1100_4/B[10] ), .Y(n2321) );
  OR2X2 U2867 ( .A(n2469), .B(\lt_x_1100_4/B[9] ), .Y(n2322) );
  AND2X2 U2868 ( .A(\lt_x_1100_4/B[8] ), .B(\sub_x_1100_2/A[8] ), .Y(n2324) );
  OR2X2 U2869 ( .A(aluOperand1[5]), .B(\lt_x_1100_4/B[5] ), .Y(n2325) );
  OR2X2 U2870 ( .A(\ashr_1100_6/SH[2] ), .B(\sub_x_1100_2/A[2] ), .Y(n2326) );
  OR2X2 U2871 ( .A(n2258), .B(aluOperand1[1]), .Y(n2327) );
  OR2X2 U2872 ( .A(\sub_x_1100_2/A[14] ), .B(n3250), .Y(n2330) );
  OR2X2 U2873 ( .A(\sub_x_1100_2/A[12] ), .B(n3251), .Y(n2331) );
  AND2X2 U2874 ( .A(n2452), .B(n3308), .Y(n2333) );
  AND2X2 U2875 ( .A(n3315), .B(n3310), .Y(n2335) );
  OR2X2 U2876 ( .A(n2261), .B(\sub_x_1100_2/A[5] ), .Y(n2337) );
  AND2X1 U2877 ( .A(n2749), .B(n2239), .Y(n2340) );
  AND2X1 U2878 ( .A(n2750), .B(n2239), .Y(n2341) );
  AND2X1 U2879 ( .A(n2752), .B(n2239), .Y(n2342) );
  AND2X1 U2880 ( .A(n2753), .B(n2239), .Y(n2343) );
  AND2X1 U2881 ( .A(n2757), .B(n2239), .Y(n2345) );
  AND2X1 U2882 ( .A(n2758), .B(n2239), .Y(n2346) );
  AND2X1 U2883 ( .A(n2759), .B(n2239), .Y(n2347) );
  AND2X2 U2884 ( .A(opcode[5]), .B(n2407), .Y(n2349) );
  INVX1 U2885 ( .A(n2351), .Y(n2352) );
  AND2X2 U2886 ( .A(n1851), .B(n4145), .Y(n2353) );
  INVX1 U2887 ( .A(n2353), .Y(n2354) );
  OR2X2 U2888 ( .A(n3725), .B(n3675), .Y(n2356) );
  AND2X2 U2889 ( .A(n1834), .B(n2268), .Y(n2357) );
  INVX1 U2890 ( .A(n2357), .Y(n2358) );
  AND2X2 U2891 ( .A(n2387), .B(n2358), .Y(n2359) );
  OR2X2 U2892 ( .A(funct3[2]), .B(\funct3[0] ), .Y(n2363) );
  OR2X2 U2893 ( .A(n3653), .B(n3726), .Y(n2364) );
  INVX1 U2894 ( .A(n2364), .Y(n2365) );
  AND2X2 U2895 ( .A(n2388), .B(n4142), .Y(n2366) );
  AND2X1 U2896 ( .A(\arithmetic_logic_unit/N149 ), .B(n4027), .Y(n2370) );
  INVX1 U2897 ( .A(n2370), .Y(n2371) );
  INVX1 U2898 ( .A(n2372), .Y(n2373) );
  INVX1 U2899 ( .A(n2374), .Y(n2375) );
  INVX1 U2900 ( .A(n2376), .Y(n2377) );
  BUFX2 U2901 ( .A(n4106), .Y(n2378) );
  BUFX2 U2902 ( .A(n4061), .Y(n2380) );
  BUFX2 U2903 ( .A(n4069), .Y(n2381) );
  OR2X2 U2904 ( .A(n3703), .B(n3702), .Y(n2382) );
  INVX1 U2905 ( .A(n2382), .Y(n2383) );
  AND2X1 U2906 ( .A(n2751), .B(n2239), .Y(n2384) );
  INVX1 U2907 ( .A(n2384), .Y(n2385) );
  AND2X2 U2908 ( .A(n1844), .B(n4168), .Y(n2386) );
  INVX1 U2909 ( .A(n2386), .Y(n2387) );
  BUFX2 U2910 ( .A(n4143), .Y(n2388) );
  BUFX2 U2911 ( .A(n4210), .Y(n2389) );
  INVX1 U2912 ( .A(n2391), .Y(n2392) );
  INVX1 U2913 ( .A(n2393), .Y(n2394) );
  AND2X2 U2914 ( .A(n3306), .B(n3314), .Y(n2395) );
  INVX1 U2915 ( .A(n2395), .Y(n2396) );
  AND2X1 U2916 ( .A(\arithmetic_logic_unit/N122 ), .B(n4027), .Y(n2397) );
  INVX1 U2917 ( .A(n2397), .Y(n2398) );
  AND2X1 U2918 ( .A(\arithmetic_logic_unit/N124 ), .B(n4027), .Y(n2399) );
  INVX1 U2919 ( .A(n2399), .Y(n2400) );
  AND2X2 U2920 ( .A(n2354), .B(n2378), .Y(n2401) );
  INVX1 U2921 ( .A(n2401), .Y(n2402) );
  AND2X2 U2922 ( .A(opcode[5]), .B(n4147), .Y(n2403) );
  INVX1 U2923 ( .A(n2403), .Y(n2404) );
  OR2X2 U2924 ( .A(opcode[3]), .B(opcode[6]), .Y(n2405) );
  INVX1 U2925 ( .A(n2405), .Y(n2406) );
  INVX1 U2926 ( .A(n2405), .Y(n2407) );
  OR2X2 U2927 ( .A(n3176), .B(n2436), .Y(n2408) );
  OR2X2 U2928 ( .A(n2438), .B(n2323), .Y(n2409) );
  INVX1 U2929 ( .A(n2409), .Y(n2410) );
  INVX1 U2930 ( .A(n2409), .Y(n2411) );
  AND2X2 U2931 ( .A(n4105), .B(opcode[4]), .Y(n2412) );
  INVX1 U2932 ( .A(n2412), .Y(n2413) );
  BUFX2 U2933 ( .A(\sub_x_1100_2/n72 ), .Y(n2414) );
  BUFX2 U2934 ( .A(\sub_x_1100_2/n90 ), .Y(n2415) );
  OR2X1 U2935 ( .A(aluOperand1[25]), .B(\lt_x_1100_4/B[25] ), .Y(n2416) );
  INVX1 U2936 ( .A(n2416), .Y(n2417) );
  OR2X1 U2937 ( .A(aluOperand1[23]), .B(\lt_x_1100_4/B[23] ), .Y(n2418) );
  INVX1 U2938 ( .A(n2418), .Y(n2419) );
  OR2X1 U2939 ( .A(aluOperand1[21]), .B(\lt_x_1100_4/B[21] ), .Y(n2420) );
  INVX1 U2940 ( .A(n2420), .Y(n2421) );
  AND2X2 U2941 ( .A(n2290), .B(n1851), .Y(n2424) );
  BUFX2 U2942 ( .A(\add_x_1100_1/n68 ), .Y(n2427) );
  BUFX2 U2943 ( .A(\add_x_1100_1/n86 ), .Y(n2428) );
  AND2X2 U2944 ( .A(n1812), .B(n2287), .Y(n2429) );
  INVX1 U2945 ( .A(n2429), .Y(n2430) );
  AND2X1 U2946 ( .A(aluOperation[0]), .B(n4103), .Y(n2431) );
  INVX1 U2947 ( .A(n2431), .Y(n2432) );
  AND2X1 U2948 ( .A(n3173), .B(n3683), .Y(n2433) );
  INVX1 U2949 ( .A(n2433), .Y(n2434) );
  AND2X2 U2950 ( .A(n2794), .B(n4322), .Y(n2435) );
  INVX1 U2951 ( .A(n2435), .Y(n2436) );
  OAI21X1 U2952 ( .A(n2882), .B(n3287), .C(n2687), .Y(n2439) );
  OR2X1 U2953 ( .A(n2236), .B(n3333), .Y(n2440) );
  INVX1 U2954 ( .A(n2440), .Y(n2441) );
  OR2X1 U2955 ( .A(n2236), .B(n3334), .Y(n2442) );
  INVX1 U2956 ( .A(n2442), .Y(n2443) );
  OR2X1 U2957 ( .A(n2236), .B(n3335), .Y(n2444) );
  INVX1 U2958 ( .A(n2444), .Y(n2445) );
  BUFX4 U2959 ( .A(aluOperand1[6]), .Y(\sub_x_1100_2/A[6] ) );
  INVX1 U2960 ( .A(n4101), .Y(n2447) );
  INVX1 U2961 ( .A(n2447), .Y(n2448) );
  INVX1 U2962 ( .A(n2450), .Y(n2449) );
  INVX1 U2963 ( .A(n2451), .Y(n2452) );
  INVX1 U2964 ( .A(n2321), .Y(n2453) );
  INVX1 U2965 ( .A(n1828), .Y(n2454) );
  INVX1 U2966 ( .A(n2454), .Y(n2455) );
  INVX1 U2967 ( .A(\add_x_1100_1/n115 ), .Y(n2456) );
  INVX1 U2968 ( .A(n2456), .Y(n2457) );
  INVX1 U2969 ( .A(\sub_x_1100_2/n119 ), .Y(n2458) );
  INVX1 U2970 ( .A(n2458), .Y(n2459) );
  BUFX2 U2971 ( .A(n2415), .Y(n2460) );
  INVX1 U2972 ( .A(n2324), .Y(n2463) );
  AND2X1 U2973 ( .A(n2793), .B(n4330), .Y(n2464) );
  INVX1 U2974 ( .A(n2464), .Y(n2465) );
  INVX1 U2975 ( .A(n2466), .Y(n2467) );
  INVX1 U2976 ( .A(n1853), .Y(n2468) );
  INVX1 U2977 ( .A(n2468), .Y(n2470) );
  OR2X1 U2978 ( .A(n3044), .B(n2472), .Y(n2471) );
  OR2X1 U2979 ( .A(n2488), .B(n2487), .Y(n2472) );
  OR2X1 U2980 ( .A(n3077), .B(n2474), .Y(n2473) );
  OR2X1 U2981 ( .A(n3075), .B(n3076), .Y(n2474) );
  OR2X1 U2982 ( .A(n3558), .B(n2476), .Y(n2475) );
  OR2X1 U2983 ( .A(n3509), .B(n3674), .Y(n2476) );
  OR2X1 U2984 ( .A(n3510), .B(n2478), .Y(n2477) );
  OR2X1 U2985 ( .A(n2490), .B(n2489), .Y(n2478) );
  AND2X2 U2986 ( .A(\sub_x_1100_2/A[2] ), .B(\ashr_1100_6/SH[2] ), .Y(n2483)
         );
  AND2X2 U2987 ( .A(aluOperand1[1]), .B(n2258), .Y(n2484) );
  OR2X1 U2988 ( .A(aluOperand1[17]), .B(n2257), .Y(n2485) );
  AND2X2 U2989 ( .A(n3725), .B(n4366), .Y(n2486) );
  OR2X1 U2990 ( .A(n4337), .B(n3304), .Y(n2487) );
  AND2X1 U2991 ( .A(\sub_x_1100_2/A[29] ), .B(n3650), .Y(n2496) );
  INVX1 U2992 ( .A(n2499), .Y(n2498) );
  AND2X1 U2993 ( .A(\arithmetic_logic_unit/N94 ), .B(n4026), .Y(n2499) );
  INVX1 U2994 ( .A(n2501), .Y(n2500) );
  AND2X1 U2995 ( .A(\arithmetic_logic_unit/N95 ), .B(n4026), .Y(n2501) );
  INVX1 U2996 ( .A(n2503), .Y(n2502) );
  INVX1 U2997 ( .A(n2505), .Y(n2504) );
  AND2X1 U2998 ( .A(n2761), .B(n2711), .Y(n2505) );
  INVX1 U2999 ( .A(n2507), .Y(n2506) );
  AND2X1 U3000 ( .A(n2762), .B(n2712), .Y(n2507) );
  INVX1 U3001 ( .A(n2509), .Y(n2508) );
  AND2X1 U3002 ( .A(n2763), .B(n2713), .Y(n2509) );
  INVX1 U3003 ( .A(n2511), .Y(n2510) );
  AND2X1 U3004 ( .A(n2764), .B(n2714), .Y(n2511) );
  INVX1 U3005 ( .A(n2513), .Y(n2512) );
  AND2X1 U3006 ( .A(n2765), .B(n2715), .Y(n2513) );
  INVX1 U3007 ( .A(n2515), .Y(n2514) );
  AND2X1 U3008 ( .A(n2766), .B(n2716), .Y(n2515) );
  INVX1 U3009 ( .A(n2517), .Y(n2516) );
  AND2X1 U3010 ( .A(n2767), .B(n2717), .Y(n2517) );
  INVX1 U3011 ( .A(n2519), .Y(n2518) );
  AND2X1 U3012 ( .A(n2768), .B(n2718), .Y(n2519) );
  INVX1 U3013 ( .A(n2521), .Y(n2520) );
  AND2X1 U3014 ( .A(n2769), .B(n2719), .Y(n2521) );
  INVX1 U3015 ( .A(n2523), .Y(n2522) );
  AND2X1 U3016 ( .A(n2770), .B(n2720), .Y(n2523) );
  INVX1 U3017 ( .A(n2525), .Y(n2524) );
  AND2X1 U3018 ( .A(n2771), .B(n2721), .Y(n2525) );
  INVX1 U3019 ( .A(n2527), .Y(n2526) );
  AND2X1 U3020 ( .A(n2772), .B(n2722), .Y(n2527) );
  INVX1 U3021 ( .A(n2529), .Y(n2528) );
  AND2X1 U3022 ( .A(n2773), .B(n2723), .Y(n2529) );
  INVX1 U3023 ( .A(n2531), .Y(n2530) );
  AND2X1 U3024 ( .A(n2774), .B(n2724), .Y(n2531) );
  INVX1 U3025 ( .A(n2533), .Y(n2532) );
  AND2X1 U3026 ( .A(n2775), .B(n2725), .Y(n2533) );
  INVX1 U3027 ( .A(n2535), .Y(n2534) );
  AND2X1 U3028 ( .A(n2776), .B(n2726), .Y(n2535) );
  INVX1 U3029 ( .A(n2537), .Y(n2536) );
  AND2X1 U3030 ( .A(n2777), .B(n2727), .Y(n2537) );
  INVX1 U3031 ( .A(n2539), .Y(n2538) );
  AND2X1 U3032 ( .A(n2778), .B(n2728), .Y(n2539) );
  INVX1 U3033 ( .A(n2541), .Y(n2540) );
  AND2X1 U3034 ( .A(n2779), .B(n2729), .Y(n2541) );
  INVX1 U3035 ( .A(n2543), .Y(n2542) );
  AND2X1 U3036 ( .A(n2780), .B(n2730), .Y(n2543) );
  INVX1 U3037 ( .A(n2545), .Y(n2544) );
  AND2X1 U3038 ( .A(n2781), .B(n2731), .Y(n2545) );
  INVX1 U3039 ( .A(n2547), .Y(n2546) );
  AND2X1 U3040 ( .A(n2782), .B(n2732), .Y(n2547) );
  INVX1 U3041 ( .A(n2549), .Y(n2548) );
  AND2X1 U3042 ( .A(n2783), .B(n2733), .Y(n2549) );
  INVX1 U3043 ( .A(n2551), .Y(n2550) );
  AND2X1 U3044 ( .A(n2784), .B(n2734), .Y(n2551) );
  INVX1 U3045 ( .A(n2553), .Y(n2552) );
  AND2X1 U3046 ( .A(n2785), .B(n2735), .Y(n2553) );
  INVX1 U3047 ( .A(n2555), .Y(n2554) );
  AND2X1 U3048 ( .A(n2786), .B(n2736), .Y(n2555) );
  INVX1 U3049 ( .A(n2557), .Y(n2556) );
  AND2X1 U3050 ( .A(n2787), .B(n2737), .Y(n2557) );
  INVX1 U3051 ( .A(n2559), .Y(n2558) );
  AND2X1 U3052 ( .A(n2788), .B(n2738), .Y(n2559) );
  INVX1 U3053 ( .A(n2561), .Y(n2560) );
  AND2X1 U3054 ( .A(n2789), .B(n2739), .Y(n2561) );
  INVX1 U3055 ( .A(n2563), .Y(n2562) );
  AND2X1 U3056 ( .A(n2790), .B(n2740), .Y(n2563) );
  INVX1 U3057 ( .A(n2565), .Y(n2564) );
  AND2X1 U3058 ( .A(n2791), .B(n2741), .Y(n2565) );
  INVX1 U3059 ( .A(n2567), .Y(n2566) );
  AND2X1 U3060 ( .A(n2792), .B(n2742), .Y(n2567) );
  INVX1 U3061 ( .A(n2569), .Y(n2568) );
  AND2X1 U3062 ( .A(n1247), .B(n3628), .Y(n2569) );
  INVX1 U3063 ( .A(n2571), .Y(n2570) );
  AND2X1 U3064 ( .A(n1247), .B(n3626), .Y(n2571) );
  INVX1 U3065 ( .A(n2573), .Y(n2572) );
  AND2X1 U3066 ( .A(n1247), .B(n3624), .Y(n2573) );
  INVX1 U3067 ( .A(n2575), .Y(n2574) );
  AND2X1 U3068 ( .A(n1247), .B(n3622), .Y(n2575) );
  INVX1 U3069 ( .A(n2577), .Y(n2576) );
  AND2X1 U3070 ( .A(n1247), .B(n3620), .Y(n2577) );
  INVX1 U3071 ( .A(n2579), .Y(n2578) );
  AND2X1 U3072 ( .A(n1247), .B(n3618), .Y(n2579) );
  INVX1 U3073 ( .A(n2581), .Y(n2580) );
  AND2X1 U3074 ( .A(n1247), .B(n3616), .Y(n2581) );
  INVX1 U3075 ( .A(n2583), .Y(n2582) );
  AND2X1 U3076 ( .A(n1247), .B(n3614), .Y(n2583) );
  INVX1 U3077 ( .A(n2585), .Y(n2584) );
  AND2X1 U3078 ( .A(n1247), .B(n3612), .Y(n2585) );
  INVX1 U3079 ( .A(n2587), .Y(n2586) );
  AND2X1 U3080 ( .A(n1247), .B(n3610), .Y(n2587) );
  INVX1 U3081 ( .A(n2589), .Y(n2588) );
  AND2X1 U3082 ( .A(n1247), .B(n3608), .Y(n2589) );
  INVX1 U3083 ( .A(n2591), .Y(n2590) );
  AND2X1 U3084 ( .A(n1247), .B(n3606), .Y(n2591) );
  INVX1 U3085 ( .A(n2593), .Y(n2592) );
  AND2X1 U3086 ( .A(n1247), .B(n3604), .Y(n2593) );
  INVX1 U3087 ( .A(n2595), .Y(n2594) );
  AND2X1 U3088 ( .A(n1247), .B(n3602), .Y(n2595) );
  INVX1 U3089 ( .A(n2597), .Y(n2596) );
  AND2X1 U3090 ( .A(n1247), .B(n3600), .Y(n2597) );
  INVX1 U3091 ( .A(n2599), .Y(n2598) );
  AND2X1 U3092 ( .A(n1247), .B(n3598), .Y(n2599) );
  INVX1 U3093 ( .A(n2601), .Y(n2600) );
  AND2X1 U3094 ( .A(n1247), .B(n3596), .Y(n2601) );
  INVX1 U3095 ( .A(n2603), .Y(n2602) );
  AND2X1 U3096 ( .A(n1247), .B(n3594), .Y(n2603) );
  INVX1 U3097 ( .A(n2605), .Y(n2604) );
  AND2X1 U3098 ( .A(n1247), .B(n3592), .Y(n2605) );
  INVX1 U3099 ( .A(n2607), .Y(n2606) );
  AND2X1 U3100 ( .A(n1247), .B(n3590), .Y(n2607) );
  INVX1 U3101 ( .A(n2609), .Y(n2608) );
  AND2X1 U3102 ( .A(n1247), .B(n3588), .Y(n2609) );
  INVX1 U3103 ( .A(n2611), .Y(n2610) );
  AND2X1 U3104 ( .A(n1247), .B(n3586), .Y(n2611) );
  INVX1 U3105 ( .A(n2613), .Y(n2612) );
  AND2X1 U3106 ( .A(n1247), .B(n3584), .Y(n2613) );
  INVX1 U3107 ( .A(n2615), .Y(n2614) );
  AND2X1 U3108 ( .A(n1247), .B(n3582), .Y(n2615) );
  INVX1 U3109 ( .A(n2617), .Y(n2616) );
  AND2X1 U3110 ( .A(n1247), .B(n3580), .Y(n2617) );
  INVX1 U3111 ( .A(n2619), .Y(n2618) );
  AND2X1 U3112 ( .A(n1247), .B(n3578), .Y(n2619) );
  INVX1 U3113 ( .A(n2621), .Y(n2620) );
  AND2X1 U3114 ( .A(n1247), .B(n3576), .Y(n2621) );
  INVX1 U3115 ( .A(n2623), .Y(n2622) );
  AND2X1 U3116 ( .A(n1247), .B(n3574), .Y(n2623) );
  INVX1 U3117 ( .A(n2625), .Y(n2624) );
  AND2X1 U3118 ( .A(n1247), .B(n3572), .Y(n2625) );
  INVX1 U3119 ( .A(n2627), .Y(n2626) );
  AND2X1 U3120 ( .A(n1247), .B(n3570), .Y(n2627) );
  INVX1 U3121 ( .A(n2629), .Y(n2628) );
  AND2X1 U3122 ( .A(n1247), .B(n3568), .Y(n2629) );
  INVX1 U3123 ( .A(n2631), .Y(n2630) );
  AND2X1 U3124 ( .A(n1247), .B(n3566), .Y(n2631) );
  AND2X2 U3125 ( .A(n4102), .B(immediate[3]), .Y(n2640) );
  INVX1 U3126 ( .A(n2640), .Y(n2641) );
  INVX1 U3127 ( .A(n2643), .Y(n2642) );
  INVX1 U3128 ( .A(n2644), .Y(n2645) );
  INVX1 U3129 ( .A(n2646), .Y(n2647) );
  INVX1 U3130 ( .A(n2649), .Y(n2648) );
  AND2X1 U3131 ( .A(n1138), .B(n4161), .Y(n2649) );
  BUFX2 U3132 ( .A(n3727), .Y(n2650) );
  BUFX2 U3133 ( .A(n3732), .Y(n2651) );
  BUFX2 U3134 ( .A(n4055), .Y(n2661) );
  INVX1 U3135 ( .A(n4059), .Y(n2663) );
  INVX1 U3136 ( .A(n2663), .Y(n2664) );
  INVX1 U3137 ( .A(n4063), .Y(n2665) );
  INVX1 U3138 ( .A(n2665), .Y(n2666) );
  INVX1 U3139 ( .A(n4065), .Y(n2667) );
  INVX1 U3140 ( .A(n2667), .Y(n2668) );
  BUFX2 U3141 ( .A(n4067), .Y(n2669) );
  BUFX2 U3142 ( .A(n4073), .Y(n2670) );
  INVX1 U3143 ( .A(n4075), .Y(n2671) );
  INVX1 U3144 ( .A(n2671), .Y(n2672) );
  INVX1 U3145 ( .A(n4077), .Y(n2673) );
  INVX1 U3146 ( .A(n2673), .Y(n2674) );
  BUFX2 U3147 ( .A(n4079), .Y(n2675) );
  INVX1 U3148 ( .A(n4081), .Y(n2676) );
  INVX1 U3149 ( .A(n2676), .Y(n2677) );
  BUFX2 U3150 ( .A(n4083), .Y(n2678) );
  BUFX2 U3151 ( .A(n4085), .Y(n2679) );
  BUFX2 U3152 ( .A(n4087), .Y(n2680) );
  BUFX2 U3153 ( .A(\add_x_1100_1/n90 ), .Y(n2682) );
  INVX1 U3154 ( .A(\add_x_1100_1/n138 ), .Y(n2683) );
  INVX1 U3155 ( .A(n2683), .Y(n2684) );
  BUFX2 U3156 ( .A(\sub_x_1100_2/n142 ), .Y(n2687) );
  AND2X1 U3157 ( .A(\sub_x_1100_2/A[27] ), .B(n3258), .Y(n2688) );
  AND2X1 U3158 ( .A(\lt_x_1100_4/B[20] ), .B(n2744), .Y(n2691) );
  INVX1 U3159 ( .A(n2339), .Y(n2692) );
  INVX1 U3160 ( .A(n2340), .Y(n2693) );
  INVX1 U3161 ( .A(n2341), .Y(n2694) );
  INVX1 U3162 ( .A(n2342), .Y(n2695) );
  INVX1 U3163 ( .A(n2343), .Y(n2696) );
  INVX1 U3164 ( .A(n2698), .Y(n2697) );
  AND2X1 U3165 ( .A(n2754), .B(n2239), .Y(n2698) );
  INVX1 U3166 ( .A(n2700), .Y(n2699) );
  AND2X1 U3167 ( .A(n2755), .B(n2239), .Y(n2700) );
  INVX1 U3168 ( .A(n2345), .Y(n2701) );
  INVX1 U3169 ( .A(n2346), .Y(n2702) );
  INVX1 U3170 ( .A(n2347), .Y(n2703) );
  INVX1 U3171 ( .A(n2348), .Y(n2704) );
  INVX1 U3172 ( .A(n2706), .Y(n2705) );
  AND2X1 U3173 ( .A(\sub_x_1100_2/A[27] ), .B(n4277), .Y(n2706) );
  INVX1 U3174 ( .A(n2708), .Y(n2707) );
  AND2X1 U3175 ( .A(\sub_x_1100_2/A[28] ), .B(n4284), .Y(n2708) );
  INVX1 U3176 ( .A(n2710), .Y(n2709) );
  AND2X2 U3177 ( .A(n1844), .B(n2223), .Y(n2710) );
  INVX1 U3178 ( .A(n2344), .Y(n2745) );
  BUFX2 U3179 ( .A(n3728), .Y(n2747) );
  INVX1 U3180 ( .A(n2356), .Y(n2794) );
  INVX1 U3181 ( .A(n2312), .Y(n2797) );
  BUFX2 U3182 ( .A(n4203), .Y(n2798) );
  BUFX2 U3183 ( .A(n4126), .Y(n2799) );
  INVX1 U3184 ( .A(n4220), .Y(n2805) );
  INVX1 U3185 ( .A(n4289), .Y(n2814) );
  INVX1 U3186 ( .A(n2814), .Y(n2815) );
  INVX1 U3187 ( .A(n2817), .Y(n2816) );
  INVX1 U3188 ( .A(n2819), .Y(n2818) );
  INVX1 U3189 ( .A(n2821), .Y(n2820) );
  INVX1 U3190 ( .A(n2823), .Y(n2822) );
  INVX1 U3191 ( .A(n2825), .Y(n2824) );
  INVX1 U3192 ( .A(n2827), .Y(n2826) );
  AND2X1 U3193 ( .A(aluOperand1[24]), .B(n3242), .Y(n2841) );
  INVX1 U3194 ( .A(n2843), .Y(n2842) );
  AND2X1 U3195 ( .A(RS1[31]), .B(n2266), .Y(n2843) );
  INVX1 U3196 ( .A(n2845), .Y(n2844) );
  AND2X1 U3197 ( .A(RS1[30]), .B(n2266), .Y(n2845) );
  INVX1 U3198 ( .A(n2847), .Y(n2846) );
  AND2X1 U3199 ( .A(RS1[29]), .B(n2266), .Y(n2847) );
  INVX1 U3200 ( .A(n2849), .Y(n2848) );
  AND2X1 U3201 ( .A(RS1[28]), .B(n2266), .Y(n2849) );
  INVX1 U3202 ( .A(n2851), .Y(n2850) );
  AND2X1 U3203 ( .A(RS1[27]), .B(n2266), .Y(n2851) );
  INVX1 U3204 ( .A(n2853), .Y(n2852) );
  AND2X1 U3205 ( .A(n3303), .B(n1144), .Y(n2853) );
  BUFX2 U3206 ( .A(n4138), .Y(n2854) );
  INVX1 U3207 ( .A(n2859), .Y(n2858) );
  AND2X1 U3208 ( .A(n3325), .B(n3781), .Y(n2859) );
  INVX1 U3209 ( .A(n2861), .Y(n2860) );
  OR2X1 U3210 ( .A(n2236), .B(n4011), .Y(n2861) );
  INVX1 U3211 ( .A(n2863), .Y(n2862) );
  OR2X1 U3212 ( .A(n2236), .B(n4014), .Y(n2863) );
  INVX1 U3213 ( .A(n2865), .Y(n2864) );
  OR2X1 U3214 ( .A(n2236), .B(n3348), .Y(n2865) );
  INVX1 U3215 ( .A(n2867), .Y(n2866) );
  INVX1 U3216 ( .A(n2869), .Y(n2868) );
  OR2X1 U3217 ( .A(n2236), .B(n3336), .Y(n2869) );
  BUFX2 U3218 ( .A(n3734), .Y(n2870) );
  OR2X2 U3219 ( .A(n3537), .B(n2797), .Y(n2871) );
  INVX1 U3220 ( .A(n2871), .Y(n2872) );
  OR2X1 U3221 ( .A(n3529), .B(n3667), .Y(n2873) );
  INVX1 U3222 ( .A(n2873), .Y(n2874) );
  BUFX2 U3223 ( .A(n3733), .Y(n2875) );
  BUFX2 U3224 ( .A(n3739), .Y(n2876) );
  BUFX2 U3225 ( .A(n3746), .Y(n2877) );
  BUFX2 U3226 ( .A(n3772), .Y(n2878) );
  INVX1 U3227 ( .A(n2881), .Y(n2880) );
  AND2X1 U3228 ( .A(n3692), .B(n2485), .Y(n2881) );
  INVX1 U3229 ( .A(n2335), .Y(n2882) );
  INVX1 U3230 ( .A(n2884), .Y(n2883) );
  AND2X1 U3231 ( .A(n4365), .B(n3553), .Y(n2884) );
  INVX1 U3232 ( .A(n2886), .Y(n2885) );
  INVX1 U3233 ( .A(n2888), .Y(n2887) );
  AND2X2 U3234 ( .A(n1145), .B(n4117), .Y(n2888) );
  BUFX2 U3235 ( .A(n3787), .Y(n2897) );
  INVX1 U3236 ( .A(n2902), .Y(n2901) );
  OR2X1 U3237 ( .A(n3907), .B(n3895), .Y(n2902) );
  INVX1 U3238 ( .A(n2904), .Y(n2903) );
  OR2X1 U3239 ( .A(n3907), .B(n3896), .Y(n2904) );
  INVX1 U3240 ( .A(n2908), .Y(n2907) );
  AND2X1 U3241 ( .A(n2251), .B(n3550), .Y(n2908) );
  INVX1 U3242 ( .A(n2910), .Y(n2909) );
  AND2X1 U3243 ( .A(n4195), .B(n2240), .Y(n2910) );
  INVX1 U3244 ( .A(n2912), .Y(n2911) );
  AND2X1 U3245 ( .A(n4200), .B(n2240), .Y(n2912) );
  INVX1 U3246 ( .A(n2915), .Y(n2914) );
  AND2X1 U3247 ( .A(n4374), .B(n4119), .Y(n2915) );
  INVX1 U3248 ( .A(n4141), .Y(n2918) );
  INVX1 U3249 ( .A(n2918), .Y(n2919) );
  INVX1 U3250 ( .A(n2921), .Y(n2920) );
  INVX1 U3251 ( .A(n2926), .Y(n2924) );
  AND2X2 U3252 ( .A(n2470), .B(n2260), .Y(n2925) );
  AND2X1 U3253 ( .A(n3238), .B(n3736), .Y(n2926) );
  INVX1 U3254 ( .A(n2928), .Y(n2927) );
  INVX1 U3255 ( .A(n2930), .Y(n2929) );
  INVX1 U3256 ( .A(n2932), .Y(n2931) );
  INVX1 U3257 ( .A(n2934), .Y(n2933) );
  INVX1 U3258 ( .A(n2936), .Y(n2935) );
  AND2X1 U3259 ( .A(instructionType[1]), .B(ir_7), .Y(n2936) );
  INVX1 U3260 ( .A(n2938), .Y(n2937) );
  AND2X1 U3261 ( .A(\arithmetic_logic_unit/N294 ), .B(aluOperation[3]), .Y(
        n2938) );
  INVX1 U3262 ( .A(n2941), .Y(n2940) );
  AND2X1 U3263 ( .A(\arithmetic_logic_unit/N268 ), .B(n4293), .Y(n2941) );
  INVX1 U3264 ( .A(n2943), .Y(n2942) );
  AND2X1 U3265 ( .A(\arithmetic_logic_unit/N272 ), .B(n4293), .Y(n2943) );
  INVX1 U3266 ( .A(n2945), .Y(n2944) );
  AND2X1 U3267 ( .A(\arithmetic_logic_unit/N273 ), .B(n4293), .Y(n2945) );
  INVX1 U3268 ( .A(n2947), .Y(n2946) );
  AND2X1 U3269 ( .A(n4293), .B(\arithmetic_logic_unit/N274 ), .Y(n2947) );
  INVX1 U3270 ( .A(n2949), .Y(n2948) );
  AND2X1 U3271 ( .A(n4293), .B(\arithmetic_logic_unit/N275 ), .Y(n2949) );
  INVX1 U3272 ( .A(n2951), .Y(n2950) );
  AND2X1 U3273 ( .A(n4293), .B(\arithmetic_logic_unit/N276 ), .Y(n2951) );
  INVX1 U3274 ( .A(n2953), .Y(n2952) );
  AND2X1 U3275 ( .A(n4293), .B(\arithmetic_logic_unit/N277 ), .Y(n2953) );
  INVX1 U3276 ( .A(n2955), .Y(n2954) );
  AND2X1 U3277 ( .A(n4293), .B(\arithmetic_logic_unit/N278 ), .Y(n2955) );
  INVX1 U3278 ( .A(n2957), .Y(n2956) );
  AND2X1 U3279 ( .A(n4293), .B(\arithmetic_logic_unit/N279 ), .Y(n2957) );
  INVX1 U3280 ( .A(n2959), .Y(n2958) );
  AND2X1 U3281 ( .A(funct7[5]), .B(n4151), .Y(n2959) );
  BUFX2 U3282 ( .A(n4256), .Y(n2969) );
  AND2X2 U3283 ( .A(aluOperation[0]), .B(n1381), .Y(n3709) );
  INVX1 U3284 ( .A(n2991), .Y(n2990) );
  AND2X1 U3285 ( .A(n3718), .B(n2413), .Y(n2991) );
  INVX1 U3286 ( .A(n2995), .Y(n2994) );
  INVX1 U3287 ( .A(n2997), .Y(n2996) );
  INVX1 U3288 ( .A(n2999), .Y(n2998) );
  INVX1 U3289 ( .A(n3001), .Y(n3000) );
  INVX1 U3290 ( .A(n3003), .Y(n3002) );
  INVX1 U3291 ( .A(n3005), .Y(n3004) );
  AND2X2 U3292 ( .A(opcode[2]), .B(n2349), .Y(n3006) );
  INVX1 U3293 ( .A(n3006), .Y(n3007) );
  INVX1 U3294 ( .A(n3009), .Y(n3008) );
  AND2X1 U3295 ( .A(n4148), .B(n3560), .Y(n3009) );
  INVX1 U3296 ( .A(n3011), .Y(n3010) );
  AND2X2 U3297 ( .A(n2220), .B(n1144), .Y(n3011) );
  INVX1 U3298 ( .A(n3013), .Y(n3012) );
  INVX1 U3299 ( .A(n3015), .Y(n3014) );
  OR2X1 U3300 ( .A(n4371), .B(ir_7), .Y(n3015) );
  INVX1 U3301 ( .A(n3017), .Y(n3016) );
  INVX1 U3302 ( .A(n3019), .Y(n3018) );
  AND2X1 U3303 ( .A(\arithmetic_logic_unit/N100 ), .B(n4026), .Y(n3019) );
  AND2X1 U3304 ( .A(\arithmetic_logic_unit/N104 ), .B(n4026), .Y(n3020) );
  INVX1 U3305 ( .A(n3022), .Y(n3021) );
  AND2X1 U3306 ( .A(\arithmetic_logic_unit/N106 ), .B(n4026), .Y(n3022) );
  INVX1 U3307 ( .A(n3024), .Y(n3023) );
  AND2X1 U3308 ( .A(\arithmetic_logic_unit/N110 ), .B(n4026), .Y(n3024) );
  INVX1 U3309 ( .A(n3026), .Y(n3025) );
  AND2X1 U3310 ( .A(\arithmetic_logic_unit/N111 ), .B(n4026), .Y(n3026) );
  INVX1 U3311 ( .A(n3028), .Y(n3027) );
  AND2X1 U3312 ( .A(\arithmetic_logic_unit/N112 ), .B(n4026), .Y(n3028) );
  INVX1 U3313 ( .A(n3030), .Y(n3029) );
  AND2X1 U3314 ( .A(\arithmetic_logic_unit/N113 ), .B(n4026), .Y(n3030) );
  INVX1 U3315 ( .A(n3032), .Y(n3031) );
  AND2X1 U3316 ( .A(\arithmetic_logic_unit/N114 ), .B(n4026), .Y(n3032) );
  INVX1 U3317 ( .A(n3034), .Y(n3033) );
  AND2X1 U3318 ( .A(\arithmetic_logic_unit/N115 ), .B(n4026), .Y(n3034) );
  INVX1 U3319 ( .A(n3036), .Y(n3035) );
  AND2X1 U3320 ( .A(\arithmetic_logic_unit/N116 ), .B(n4026), .Y(n3036) );
  INVX1 U3321 ( .A(n3038), .Y(n3037) );
  AND2X1 U3322 ( .A(funct3[1]), .B(n1145), .Y(n3038) );
  INVX1 U3323 ( .A(n3041), .Y(n3040) );
  AND2X1 U3324 ( .A(memoryReady), .B(n2269), .Y(n3041) );
  INVX1 U3325 ( .A(n3043), .Y(n3042) );
  AND2X1 U3326 ( .A(n4129), .B(n3172), .Y(n3043) );
  INVX1 U3327 ( .A(n3296), .Y(n3044) );
  INVX1 U3328 ( .A(n3047), .Y(n3046) );
  AND2X2 U3329 ( .A(n2358), .B(n3296), .Y(n3047) );
  INVX1 U3330 ( .A(n3049), .Y(n3048) );
  INVX1 U3331 ( .A(n3051), .Y(n3050) );
  AND2X1 U3332 ( .A(n4367), .B(n1139), .Y(n3051) );
  INVX1 U3333 ( .A(n3053), .Y(n3052) );
  AND2X1 U3334 ( .A(n3517), .B(funct7[5]), .Y(n3053) );
  INVX1 U3335 ( .A(n3056), .Y(n3055) );
  INVX1 U3336 ( .A(n3067), .Y(n3066) );
  AND2X1 U3337 ( .A(n3212), .B(\add_x_1100_1/n197 ), .Y(n3067) );
  INVX1 U3338 ( .A(n3069), .Y(n3068) );
  AND2X1 U3339 ( .A(n3236), .B(n3289), .Y(n3069) );
  BUFX2 U3340 ( .A(n533), .Y(n3071) );
  INVX1 U3341 ( .A(n4178), .Y(n3075) );
  INVX1 U3342 ( .A(n4179), .Y(n3076) );
  INVX1 U3343 ( .A(n4180), .Y(n3077) );
  BUFX2 U3344 ( .A(n967), .Y(n3094) );
  INVX1 U3345 ( .A(n3096), .Y(n3095) );
  AND2X1 U3346 ( .A(n3723), .B(funct7[0]), .Y(n3096) );
  INVX1 U3347 ( .A(n3098), .Y(n3097) );
  AND2X1 U3348 ( .A(n3723), .B(funct7[1]), .Y(n3098) );
  INVX1 U3349 ( .A(n3100), .Y(n3099) );
  AND2X1 U3350 ( .A(n3723), .B(funct7[2]), .Y(n3100) );
  INVX1 U3351 ( .A(n3102), .Y(n3101) );
  AND2X1 U3352 ( .A(n3723), .B(funct7[3]), .Y(n3102) );
  INVX1 U3353 ( .A(n3104), .Y(n3103) );
  AND2X1 U3354 ( .A(n3723), .B(funct7[4]), .Y(n3104) );
  INVX1 U3355 ( .A(n3106), .Y(n3105) );
  AND2X1 U3356 ( .A(n3723), .B(funct7[5]), .Y(n3106) );
  INVX1 U3357 ( .A(n3109), .Y(n3108) );
  INVX1 U3358 ( .A(n3111), .Y(n3110) );
  AND2X1 U3359 ( .A(n3649), .B(n3686), .Y(n3111) );
  INVX1 U3360 ( .A(n3113), .Y(n3112) );
  AND2X1 U3361 ( .A(n2159), .B(n3688), .Y(n3113) );
  INVX1 U3362 ( .A(n3115), .Y(n3114) );
  AND2X1 U3363 ( .A(n3644), .B(n3689), .Y(n3115) );
  INVX1 U3364 ( .A(n3117), .Y(n3116) );
  AND2X1 U3365 ( .A(n2088), .B(n3690), .Y(n3117) );
  INVX1 U3366 ( .A(n3119), .Y(n3118) );
  AND2X1 U3367 ( .A(n2229), .B(n3666), .Y(n3119) );
  INVX1 U3368 ( .A(n3121), .Y(n3120) );
  AND2X1 U3369 ( .A(n3188), .B(n3259), .Y(n3121) );
  INVX1 U3370 ( .A(n3123), .Y(n3122) );
  AND2X1 U3371 ( .A(n3190), .B(n2416), .Y(n3123) );
  INVX1 U3372 ( .A(n3125), .Y(n3124) );
  AND2X1 U3373 ( .A(n3192), .B(n2418), .Y(n3125) );
  INVX1 U3374 ( .A(n3127), .Y(n3126) );
  AND2X1 U3375 ( .A(n3194), .B(n2420), .Y(n3127) );
  INVX1 U3376 ( .A(n3129), .Y(n3128) );
  AND2X1 U3377 ( .A(n3199), .B(n2313), .Y(n3129) );
  INVX1 U3378 ( .A(n3131), .Y(n3130) );
  AND2X1 U3379 ( .A(n3203), .B(\add_x_1100_1/n187 ), .Y(n3131) );
  INVX1 U3380 ( .A(n3133), .Y(n3132) );
  AND2X1 U3381 ( .A(n2482), .B(\add_x_1100_1/n192 ), .Y(n3133) );
  INVX1 U3382 ( .A(n3135), .Y(n3134) );
  AND2X1 U3383 ( .A(n3208), .B(\add_x_1100_1/n193 ), .Y(n3135) );
  INVX1 U3384 ( .A(n3137), .Y(n3136) );
  AND2X1 U3385 ( .A(n3213), .B(n3260), .Y(n3137) );
  INVX1 U3386 ( .A(n3139), .Y(n3138) );
  AND2X1 U3387 ( .A(n3215), .B(n3262), .Y(n3139) );
  INVX1 U3388 ( .A(n3141), .Y(n3140) );
  AND2X1 U3389 ( .A(n3217), .B(n3263), .Y(n3141) );
  INVX1 U3390 ( .A(n3143), .Y(n3142) );
  AND2X1 U3391 ( .A(n3219), .B(n3265), .Y(n3143) );
  INVX1 U3392 ( .A(n3145), .Y(n3144) );
  AND2X1 U3393 ( .A(n3640), .B(n2485), .Y(n3145) );
  INVX1 U3394 ( .A(n3147), .Y(n3146) );
  AND2X1 U3395 ( .A(n3223), .B(n3659), .Y(n3147) );
  INVX1 U3396 ( .A(n3149), .Y(n3148) );
  AND2X1 U3397 ( .A(n3227), .B(n2334), .Y(n3149) );
  INVX1 U3398 ( .A(n3151), .Y(n3150) );
  AND2X1 U3399 ( .A(n3669), .B(n3539), .Y(n3151) );
  INVX1 U3400 ( .A(n3153), .Y(n3152) );
  AND2X1 U3401 ( .A(n3233), .B(\sub_x_1100_2/n198 ), .Y(n3153) );
  INVX1 U3402 ( .A(n3155), .Y(n3154) );
  AND2X1 U3403 ( .A(\lt_x_1100_4/B[26] ), .B(aluOperand1[26]), .Y(n3156) );
  INVX1 U3404 ( .A(n3158), .Y(n3157) );
  AND2X1 U3405 ( .A(\lt_x_1100_4/B[24] ), .B(aluOperand1[24]), .Y(n3158) );
  AND2X1 U3406 ( .A(\lt_x_1100_4/B[22] ), .B(aluOperand1[22]), .Y(n3159) );
  AND2X1 U3407 ( .A(\lt_x_1100_4/B[20] ), .B(aluOperand1[20]), .Y(n3160) );
  AND2X1 U3408 ( .A(\sub_x_1100_2/n216 ), .B(aluOperand1[18]), .Y(n3162) );
  INVX1 U3409 ( .A(n3163), .Y(n3164) );
  INVX1 U3410 ( .A(n3166), .Y(n3165) );
  AND2X2 U3411 ( .A(n2221), .B(n2406), .Y(n3167) );
  INVX1 U3412 ( .A(n3172), .Y(n3171) );
  OR2X2 U3413 ( .A(n3562), .B(n2437), .Y(n3172) );
  INVX1 U3414 ( .A(n3174), .Y(n3173) );
  INVX1 U3415 ( .A(n2355), .Y(n3176) );
  INVX1 U3416 ( .A(n2446), .Y(n3181) );
  INVX1 U3417 ( .A(n2314), .Y(n3182) );
  INVX1 U3418 ( .A(n2315), .Y(n3185) );
  AND2X2 U3419 ( .A(n3726), .B(n4130), .Y(n3186) );
  INVX1 U3420 ( .A(n3189), .Y(n3188) );
  AND2X1 U3421 ( .A(\lt_x_1100_4/B[27] ), .B(\sub_x_1100_2/A[27] ), .Y(n3189)
         );
  INVX1 U3422 ( .A(n3191), .Y(n3190) );
  AND2X1 U3423 ( .A(\lt_x_1100_4/B[25] ), .B(aluOperand1[25]), .Y(n3191) );
  INVX1 U3424 ( .A(n3193), .Y(n3192) );
  AND2X1 U3425 ( .A(\lt_x_1100_4/B[23] ), .B(aluOperand1[23]), .Y(n3193) );
  INVX1 U3426 ( .A(n3195), .Y(n3194) );
  AND2X1 U3427 ( .A(\lt_x_1100_4/B[21] ), .B(aluOperand1[21]), .Y(n3195) );
  INVX1 U3428 ( .A(n3197), .Y(n3196) );
  AND2X1 U3429 ( .A(\lt_x_1100_4/B[19] ), .B(aluOperand1[19]), .Y(n3197) );
  INVX1 U3430 ( .A(n3207), .Y(n3206) );
  INVX1 U3431 ( .A(n3209), .Y(n3208) );
  AND2X2 U3432 ( .A(aluOperand1[3]), .B(n1821), .Y(n3210) );
  INVX1 U3433 ( .A(n3210), .Y(n3211) );
  INVX1 U3434 ( .A(n2484), .Y(n3212) );
  INVX1 U3435 ( .A(n3214), .Y(n3213) );
  AND2X1 U3436 ( .A(n3258), .B(\sub_x_1100_2/A[27] ), .Y(n3214) );
  INVX1 U3437 ( .A(n3216), .Y(n3215) );
  AND2X1 U3438 ( .A(n3241), .B(aluOperand1[25]), .Y(n3216) );
  INVX1 U3439 ( .A(n3218), .Y(n3217) );
  AND2X1 U3440 ( .A(n3243), .B(aluOperand1[23]), .Y(n3218) );
  INVX1 U3441 ( .A(n3220), .Y(n3219) );
  AND2X1 U3442 ( .A(n3245), .B(aluOperand1[21]), .Y(n3220) );
  INVX1 U3443 ( .A(n3222), .Y(n3221) );
  AND2X1 U3444 ( .A(n3247), .B(aluOperand1[19]), .Y(n3222) );
  INVX1 U3445 ( .A(n3224), .Y(n3223) );
  INVX1 U3446 ( .A(n3226), .Y(n3225) );
  INVX1 U3447 ( .A(n3228), .Y(n3227) );
  INVX1 U3448 ( .A(n3230), .Y(n3229) );
  AND2X2 U3449 ( .A(n2260), .B(n2470), .Y(n3230) );
  INVX1 U3450 ( .A(n3232), .Y(n3231) );
  INVX1 U3451 ( .A(n3234), .Y(n3233) );
  INVX1 U3452 ( .A(n3237), .Y(n3236) );
  BUFX2 U3453 ( .A(n4214), .Y(n3250) );
  BUFX2 U3454 ( .A(n4212), .Y(n3251) );
  BUFX2 U3455 ( .A(n4205), .Y(n3252) );
  INVX1 U3456 ( .A(n3254), .Y(n3253) );
  AND2X1 U3457 ( .A(n2454), .B(n3321), .Y(n3254) );
  OR2X1 U3458 ( .A(\sub_x_1100_2/A[27] ), .B(\lt_x_1100_4/B[27] ), .Y(n3259)
         );
  OR2X1 U3459 ( .A(\sub_x_1100_2/A[27] ), .B(n3258), .Y(n3260) );
  INVX1 U3460 ( .A(n3262), .Y(n3261) );
  OR2X1 U3461 ( .A(aluOperand1[25]), .B(n3241), .Y(n3262) );
  OR2X1 U3462 ( .A(aluOperand1[23]), .B(n3243), .Y(n3263) );
  INVX1 U3463 ( .A(n3265), .Y(n3264) );
  OR2X1 U3464 ( .A(aluOperand1[21]), .B(n3245), .Y(n3265) );
  INVX1 U3465 ( .A(n3267), .Y(n3266) );
  OR2X1 U3466 ( .A(aluOperand1[19]), .B(n3247), .Y(n3267) );
  INVX1 U3467 ( .A(n3278), .Y(n3277) );
  BUFX2 U3468 ( .A(n3955), .Y(n3278) );
  BUFX2 U3469 ( .A(n3967), .Y(n3279) );
  BUFX2 U3470 ( .A(n2428), .Y(n3284) );
  INVX1 U3471 ( .A(\add_x_1100_1/n157 ), .Y(n3285) );
  INVX1 U3472 ( .A(n3285), .Y(n3286) );
  BUFX2 U3473 ( .A(\sub_x_1100_2/n161 ), .Y(n3287) );
  INVX1 U3474 ( .A(n3291), .Y(n3290) );
  OR2X1 U3475 ( .A(n2238), .B(n3364), .Y(n3291) );
  INVX1 U3476 ( .A(n3293), .Y(n3292) );
  OR2X1 U3477 ( .A(n2238), .B(n3939), .Y(n3293) );
  INVX1 U3478 ( .A(n3295), .Y(n3294) );
  OR2X1 U3479 ( .A(n2238), .B(n3365), .Y(n3295) );
  INVX1 U3480 ( .A(n3297), .Y(n3298) );
  OR2X2 U3481 ( .A(n1145), .B(n2220), .Y(n3302) );
  OR2X2 U3482 ( .A(n3178), .B(n3540), .Y(n3305) );
  INVX1 U3483 ( .A(n3305), .Y(n3306) );
  INVX1 U3484 ( .A(n3307), .Y(n3308) );
  OR2X2 U3485 ( .A(n3180), .B(n2338), .Y(n3309) );
  INVX1 U3486 ( .A(n3309), .Y(n3310) );
  INVX1 U3487 ( .A(n3312), .Y(n3311) );
  OR2X2 U3488 ( .A(n3181), .B(n2480), .Y(n3313) );
  INVX1 U3489 ( .A(n3313), .Y(n3314) );
  INVX1 U3490 ( .A(n3316), .Y(n3315) );
  OR2X1 U3491 ( .A(n3534), .B(n3538), .Y(n3316) );
  BUFX2 U3492 ( .A(n2457), .Y(n3317) );
  BUFX2 U3493 ( .A(n2268), .Y(n3318) );
  INVX1 U3494 ( .A(n3320), .Y(n3319) );
  AND2X2 U3495 ( .A(n3164), .B(n3298), .Y(n3320) );
  INVX1 U3496 ( .A(n3322), .Y(n3321) );
  INVX1 U3497 ( .A(n3324), .Y(n3323) );
  OR2X1 U3498 ( .A(n1841), .B(n3363), .Y(n3324) );
  BUFX2 U3499 ( .A(n3882), .Y(n3328) );
  BUFX2 U3500 ( .A(n3988), .Y(n3332) );
  INVX1 U3501 ( .A(n2333), .Y(n3337) );
  INVX1 U3502 ( .A(n3339), .Y(n3338) );
  INVX1 U3503 ( .A(n3341), .Y(n3340) );
  AND2X1 U3504 ( .A(n3858), .B(n3908), .Y(n3341) );
  INVX1 U3505 ( .A(n3343), .Y(n3342) );
  AND2X1 U3506 ( .A(n3824), .B(n3908), .Y(n3343) );
  INVX1 U3507 ( .A(n3345), .Y(n3344) );
  AND2X1 U3508 ( .A(n3828), .B(n3908), .Y(n3345) );
  INVX1 U3509 ( .A(n3346), .Y(n3347) );
  INVX1 U3510 ( .A(n3349), .Y(n3348) );
  INVX1 U3511 ( .A(n3351), .Y(n3350) );
  INVX1 U3512 ( .A(n3353), .Y(n3352) );
  AND2X1 U3513 ( .A(n3968), .B(n3908), .Y(n3353) );
  INVX1 U3514 ( .A(n3367), .Y(n3366) );
  INVX1 U3515 ( .A(n3369), .Y(n3368) );
  INVX1 U3516 ( .A(n4146), .Y(n3377) );
  INVX1 U3517 ( .A(n3377), .Y(n3378) );
  BUFX2 U3518 ( .A(n3842), .Y(n3421) );
  BUFX2 U3519 ( .A(n3880), .Y(n3423) );
  BUFX2 U3520 ( .A(n3932), .Y(n3470) );
  BUFX2 U3521 ( .A(n3931), .Y(n3471) );
  BUFX2 U3522 ( .A(n3936), .Y(n3474) );
  BUFX2 U3523 ( .A(n3996), .Y(n3489) );
  INVX1 U3524 ( .A(n3502), .Y(n3501) );
  INVX1 U3525 ( .A(n3504), .Y(n3503) );
  OR2X2 U3526 ( .A(n3724), .B(n2212), .Y(n3505) );
  INVX1 U3527 ( .A(n3508), .Y(n3507) );
  INVX1 U3528 ( .A(n2437), .Y(n3509) );
  INVX1 U3529 ( .A(n4325), .Y(n3510) );
  OR2X1 U3530 ( .A(aluOperation[1]), .B(aluOperation[2]), .Y(n245) );
  BUFX2 U3531 ( .A(n2052), .Y(n3511) );
  BUFX2 U3532 ( .A(n2051), .Y(n3512) );
  BUFX2 U3533 ( .A(n2058), .Y(n3514) );
  BUFX2 U3534 ( .A(n2059), .Y(n3515) );
  INVX1 U3535 ( .A(n3521), .Y(n3520) );
  AND2X2 U3536 ( .A(aluOperand1[4]), .B(\sub_x_1100_2/B[4] ), .Y(n3521) );
  INVX1 U3537 ( .A(n3525), .Y(n3524) );
  INVX1 U3538 ( .A(n2320), .Y(n3532) );
  INVX1 U3539 ( .A(n2336), .Y(n3534) );
  BUFX2 U3540 ( .A(n3181), .Y(n3536) );
  INVX1 U3541 ( .A(n2326), .Y(n3537) );
  INVX1 U3542 ( .A(n3539), .Y(n3538) );
  INVX1 U3543 ( .A(n2325), .Y(n3540) );
  INVX1 U3544 ( .A(n2483), .Y(n3541) );
  INVX1 U3545 ( .A(n3543), .Y(n3542) );
  AND2X2 U3546 ( .A(n2259), .B(\sub_x_1100_2/A[8] ), .Y(n3543) );
  INVX1 U3547 ( .A(n3547), .Y(n3546) );
  AND2X2 U3548 ( .A(opcode[2]), .B(n2222), .Y(n3547) );
  AND2X2 U3549 ( .A(n3562), .B(n2270), .Y(n4108) );
  INVX1 U3550 ( .A(n4140), .Y(n3551) );
  INVX1 U3551 ( .A(n3551), .Y(n3552) );
  INVX1 U3552 ( .A(n3551), .Y(n3553) );
  BUFX2 U3553 ( .A(n2288), .Y(n3555) );
  OR2X1 U3554 ( .A(funct7[6]), .B(instructionType[2]), .Y(n4181) );
  INVX1 U3555 ( .A(n2329), .Y(n3556) );
  INVX1 U3556 ( .A(n1826), .Y(n3557) );
  BUFX2 U3557 ( .A(n1103), .Y(n3559) );
  BUFX2 U3558 ( .A(n2267), .Y(n3560) );
  BUFX2 U3559 ( .A(n4317), .Y(n3563) );
  BUFX2 U3560 ( .A(n4314), .Y(n3564) );
  AND2X1 U3561 ( .A(n4030), .B(N1117), .Y(n3565) );
  INVX1 U3562 ( .A(n3565), .Y(n3566) );
  AND2X1 U3563 ( .A(n4030), .B(N1120), .Y(n3567) );
  INVX1 U3564 ( .A(n3567), .Y(n3568) );
  AND2X1 U3565 ( .A(n4030), .B(N1123), .Y(n3569) );
  INVX1 U3566 ( .A(n3569), .Y(n3570) );
  AND2X1 U3567 ( .A(n4030), .B(N1126), .Y(n3571) );
  INVX1 U3568 ( .A(n3571), .Y(n3572) );
  AND2X1 U3569 ( .A(n4030), .B(N1129), .Y(n3573) );
  INVX1 U3570 ( .A(n3573), .Y(n3574) );
  AND2X1 U3571 ( .A(n4030), .B(N1132), .Y(n3575) );
  INVX1 U3572 ( .A(n3575), .Y(n3576) );
  AND2X1 U3573 ( .A(n4030), .B(N1135), .Y(n3577) );
  INVX1 U3574 ( .A(n3577), .Y(n3578) );
  AND2X1 U3575 ( .A(n4030), .B(N1138), .Y(n3579) );
  INVX1 U3576 ( .A(n3579), .Y(n3580) );
  AND2X1 U3577 ( .A(n4030), .B(N1141), .Y(n3581) );
  INVX1 U3578 ( .A(n3581), .Y(n3582) );
  AND2X1 U3579 ( .A(n4030), .B(N1144), .Y(n3583) );
  INVX1 U3580 ( .A(n3583), .Y(n3584) );
  AND2X1 U3581 ( .A(n4030), .B(N1147), .Y(n3585) );
  INVX1 U3582 ( .A(n3585), .Y(n3586) );
  AND2X1 U3583 ( .A(n4030), .B(N1150), .Y(n3587) );
  INVX1 U3584 ( .A(n3587), .Y(n3588) );
  AND2X1 U3585 ( .A(n4030), .B(N1153), .Y(n3589) );
  INVX1 U3586 ( .A(n3589), .Y(n3590) );
  AND2X1 U3587 ( .A(n4030), .B(N1156), .Y(n3591) );
  INVX1 U3588 ( .A(n3591), .Y(n3592) );
  AND2X1 U3589 ( .A(n4030), .B(N1159), .Y(n3593) );
  INVX1 U3590 ( .A(n3593), .Y(n3594) );
  AND2X1 U3591 ( .A(n4030), .B(N1162), .Y(n3595) );
  INVX1 U3592 ( .A(n3595), .Y(n3596) );
  AND2X1 U3593 ( .A(n4030), .B(N1165), .Y(n3597) );
  INVX1 U3594 ( .A(n3597), .Y(n3598) );
  INVX1 U3595 ( .A(n3599), .Y(n3600) );
  AND2X1 U3596 ( .A(n4030), .B(N1171), .Y(n3601) );
  INVX1 U3597 ( .A(n3601), .Y(n3602) );
  INVX1 U3598 ( .A(n3603), .Y(n3604) );
  AND2X1 U3599 ( .A(n4030), .B(N1177), .Y(n3605) );
  INVX1 U3600 ( .A(n3605), .Y(n3606) );
  AND2X1 U3601 ( .A(n4030), .B(N1180), .Y(n3607) );
  INVX1 U3602 ( .A(n3607), .Y(n3608) );
  AND2X1 U3603 ( .A(n4030), .B(N1183), .Y(n3609) );
  INVX1 U3604 ( .A(n3609), .Y(n3610) );
  AND2X1 U3605 ( .A(n4030), .B(N1186), .Y(n3611) );
  INVX1 U3606 ( .A(n3611), .Y(n3612) );
  AND2X1 U3607 ( .A(n4030), .B(N1189), .Y(n3613) );
  INVX1 U3608 ( .A(n3613), .Y(n3614) );
  AND2X1 U3609 ( .A(n4030), .B(N1192), .Y(n3615) );
  INVX1 U3610 ( .A(n3615), .Y(n3616) );
  INVX1 U3611 ( .A(n3617), .Y(n3618) );
  INVX1 U3612 ( .A(n3619), .Y(n3620) );
  INVX1 U3613 ( .A(n3621), .Y(n3622) );
  INVX1 U3614 ( .A(n3623), .Y(n3624) );
  AND2X1 U3615 ( .A(n4030), .B(N1207), .Y(n3625) );
  INVX1 U3616 ( .A(n3625), .Y(n3626) );
  AND2X1 U3617 ( .A(n4030), .B(N1210), .Y(n3627) );
  INVX1 U3618 ( .A(n3627), .Y(n3628) );
  BUFX2 U3619 ( .A(n963), .Y(n3629) );
  BUFX2 U3620 ( .A(n955), .Y(n3630) );
  INVX1 U3621 ( .A(n3631), .Y(n3632) );
  AND2X1 U3622 ( .A(\opcode[1] ), .B(\opcode[0] ), .Y(n4325) );
  INVX1 U3623 ( .A(n3633), .Y(n3634) );
  INVX1 U3624 ( .A(n3635), .Y(n3636) );
  INVX1 U3625 ( .A(n3637), .Y(n3638) );
  INVX1 U3626 ( .A(n3639), .Y(n3640) );
  AND2X1 U3627 ( .A(n3240), .B(aluOperand1[26]), .Y(n3641) );
  AND2X1 U3628 ( .A(n3244), .B(aluOperand1[22]), .Y(n3642) );
  AND2X1 U3629 ( .A(n3242), .B(aluOperand1[24]), .Y(n3643) );
  INVX1 U3630 ( .A(n3643), .Y(n3644) );
  AND2X1 U3631 ( .A(n3246), .B(aluOperand1[20]), .Y(n3645) );
  AND2X1 U3632 ( .A(\lt_x_1100_4/B[18] ), .B(aluOperand1[18]), .Y(n3647) );
  AND2X1 U3633 ( .A(n3257), .B(\sub_x_1100_2/A[28] ), .Y(n3648) );
  INVX1 U3634 ( .A(n3648), .Y(n3649) );
  BUFX2 U3635 ( .A(n4290), .Y(n3650) );
  AND2X1 U3636 ( .A(n2240), .B(n2241), .Y(n3651) );
  OR2X1 U3637 ( .A(n4117), .B(aluSignRegister), .Y(n3652) );
  INVX1 U3638 ( .A(n3652), .Y(n3653) );
  BUFX2 U3639 ( .A(n3982), .Y(n3654) );
  AND2X1 U3640 ( .A(n4364), .B(pcWrite), .Y(n4340) );
  INVX1 U3641 ( .A(n3659), .Y(n3660) );
  INVX1 U3642 ( .A(n3668), .Y(n3669) );
  BUFX2 U3643 ( .A(n4194), .Y(n3670) );
  INVX1 U3644 ( .A(n3670), .Y(n3907) );
  INVX1 U3645 ( .A(memoryReadWrite), .Y(n1001) );
  OR2X2 U3646 ( .A(opcode[2]), .B(opcode[3]), .Y(n3671) );
  INVX1 U3647 ( .A(n3671), .Y(n3672) );
  BUFX2 U3648 ( .A(n987), .Y(n3675) );
  AND2X2 U3649 ( .A(n3675), .B(n3725), .Y(n4130) );
  AND2X1 U3650 ( .A(n3723), .B(n4367), .Y(n3676) );
  INVX1 U3651 ( .A(n3676), .Y(n3677) );
  INVX1 U3652 ( .A(instructionOrData), .Y(n1034) );
  OR2X1 U3653 ( .A(aluOperand1[24]), .B(\lt_x_1100_4/B[24] ), .Y(n3678) );
  OR2X1 U3654 ( .A(aluOperand1[22]), .B(\lt_x_1100_4/B[22] ), .Y(n3679) );
  OR2X1 U3655 ( .A(aluOperand1[20]), .B(\lt_x_1100_4/B[20] ), .Y(n3680) );
  OR2X1 U3656 ( .A(aluOperand1[26]), .B(\lt_x_1100_4/B[26] ), .Y(n3681) );
  OR2X1 U3657 ( .A(aluOperand1[18]), .B(\lt_x_1100_4/B[18] ), .Y(n3682) );
  OR2X1 U3658 ( .A(aluOperand1[17]), .B(\lt_x_1100_4/B[17] ), .Y(n3683) );
  OR2X1 U3659 ( .A(aluOperand1[16]), .B(\lt_x_1100_4/B[16] ), .Y(n3684) );
  INVX1 U3660 ( .A(\add_x_1100_1/n136 ), .Y(\add_x_1100_1/n135 ) );
  INVX1 U3661 ( .A(\add_x_1100_1/n166 ), .Y(\add_x_1100_1/n165 ) );
  INVX1 U3662 ( .A(n2291), .Y(\add_x_1100_1/n156 ) );
  INVX1 U3663 ( .A(n3284), .Y(\add_x_1100_1/n85 ) );
  INVX1 U3664 ( .A(n2411), .Y(\add_x_1100_1/n126 ) );
  INVX1 U3665 ( .A(\add_x_1100_1/n129 ), .Y(\add_x_1100_1/n127 ) );
  INVX1 U3666 ( .A(n2453), .Y(\add_x_1100_1/n188 ) );
  INVX1 U3667 ( .A(n2328), .Y(\add_x_1100_1/n197 ) );
  INVX1 U3668 ( .A(\add_x_1100_1/n113 ), .Y(\add_x_1100_1/n112 ) );
  INVX1 U3669 ( .A(n3185), .Y(\add_x_1100_1/n186 ) );
  INVX1 U3670 ( .A(\add_x_1100_1/n104 ), .Y(\add_x_1100_1/n102 ) );
  INVX1 U3671 ( .A(n3182), .Y(\add_x_1100_1/n96 ) );
  INVX1 U3672 ( .A(n2273), .Y(\add_x_1100_1/n193 ) );
  INVX1 U3673 ( .A(n3532), .Y(\add_x_1100_1/n187 ) );
  INVX1 U3674 ( .A(n2797), .Y(\add_x_1100_1/n195 ) );
  INVX1 U3675 ( .A(n3536), .Y(\add_x_1100_1/n192 ) );
  OR2X1 U3676 ( .A(\sub_x_1100_2/A[28] ), .B(n3257), .Y(n3686) );
  OR2X1 U3677 ( .A(aluOperand1[18]), .B(\sub_x_1100_2/n216 ), .Y(n3687) );
  OR2X1 U3678 ( .A(aluOperand1[26]), .B(n3240), .Y(n3688) );
  OR2X1 U3679 ( .A(aluOperand1[24]), .B(n3242), .Y(n3689) );
  OR2X1 U3680 ( .A(aluOperand1[22]), .B(n3244), .Y(n3690) );
  OR2X1 U3681 ( .A(aluOperand1[20]), .B(n3246), .Y(n3691) );
  OR2X1 U3682 ( .A(aluOperand1[16]), .B(n2263), .Y(n3692) );
  INVX1 U3683 ( .A(\lt_x_1100_4/B[7] ), .Y(\sub_x_1100_2/n227 ) );
  INVX1 U3684 ( .A(\lt_x_1100_4/B[6] ), .Y(\sub_x_1100_2/n228 ) );
  INVX1 U3685 ( .A(n1823), .Y(n3685) );
  INVX1 U3686 ( .A(\lt_x_1100_4/B[18] ), .Y(\sub_x_1100_2/n216 ) );
  INVX1 U3687 ( .A(n2217), .Y(\sub_x_1100_2/n139 ) );
  INVX1 U3688 ( .A(\sub_x_1100_2/n170 ), .Y(\sub_x_1100_2/n169 ) );
  INVX1 U3689 ( .A(n1822), .Y(\sub_x_1100_2/n160 ) );
  INVX1 U3690 ( .A(n2460), .Y(\sub_x_1100_2/n89 ) );
  INVX1 U3691 ( .A(\sub_x_1100_2/n133 ), .Y(\sub_x_1100_2/n131 ) );
  INVX1 U3692 ( .A(\sub_x_1100_2/n117 ), .Y(\sub_x_1100_2/n116 ) );
  INVX1 U3693 ( .A(\sub_x_1100_2/n108 ), .Y(\sub_x_1100_2/n106 ) );
  INVX1 U3694 ( .A(n2338), .Y(\sub_x_1100_2/n198 ) );
  INVX1 U3695 ( .A(n3694), .Y(n3695) );
  INVX1 U3696 ( .A(n3694), .Y(n3696) );
  INVX1 U3697 ( .A(n3693), .Y(n3697) );
  INVX1 U3698 ( .A(n3694), .Y(n3698) );
  INVX1 U3699 ( .A(n3694), .Y(n3699) );
  INVX1 U3700 ( .A(n3694), .Y(n3700) );
  INVX1 U3701 ( .A(n3694), .Y(n3701) );
  BUFX4 U3702 ( .A(aluOperand1[5]), .Y(\sub_x_1100_2/A[5] ) );
  BUFX4 U3703 ( .A(aluOperand1[2]), .Y(\sub_x_1100_2/A[2] ) );
  BUFX4 U3704 ( .A(aluOperand1[8]), .Y(\sub_x_1100_2/A[8] ) );
  INVX2 U3705 ( .A(n2437), .Y(n4168) );
  AND2X2 U3706 ( .A(n2352), .B(n2641), .Y(n3712) );
  AND2X2 U3707 ( .A(n2448), .B(n2642), .Y(n3707) );
  INVX8 U3708 ( .A(n4036), .Y(n4091) );
  INVX1 U3709 ( .A(n3715), .Y(n4028) );
  AND2X2 U3710 ( .A(n2647), .B(n2377), .Y(n3706) );
  INVX1 U3711 ( .A(n3708), .Y(n4031) );
  OR2X1 U3712 ( .A(n2828), .B(n3562), .Y(n4034) );
  AND2X1 U3713 ( .A(instructionType[2]), .B(n4370), .Y(n3717) );
  OR2X1 U3714 ( .A(n3166), .B(n245), .Y(n3711) );
  INVX1 U3715 ( .A(aluOperation[3]), .Y(n4103) );
  INVX1 U3716 ( .A(funct7[6]), .Y(n4367) );
  AND2X2 U3717 ( .A(n2645), .B(n2375), .Y(n3705) );
  AND2X1 U3718 ( .A(n4371), .B(n4370), .Y(n4173) );
  INVX1 U3719 ( .A(n3717), .Y(n3723) );
  INVX1 U3720 ( .A(instructionType[0]), .Y(n4370) );
  INVX1 U3721 ( .A(instructionType[1]), .Y(n4371) );
  INVX1 U3722 ( .A(instructionType[2]), .Y(n4372) );
  INVX1 U3723 ( .A(n3724), .Y(n4365) );
  INVX1 U3724 ( .A(n3726), .Y(n4334) );
  BUFX2 U3725 ( .A(n1000), .Y(n3726) );
  BUFX2 U3726 ( .A(n995), .Y(n3724) );
  AND2X2 U3727 ( .A(n3165), .B(n4104), .Y(n3704) );
  AND2X2 U3728 ( .A(aluSrcA[1]), .B(n4035), .Y(n4036) );
  AND2X2 U3729 ( .A(aluSrcA[0]), .B(n2274), .Y(n4089) );
  AND2X2 U3730 ( .A(aluSrcB[1]), .B(n4092), .Y(n4102) );
  INVX1 U3731 ( .A(n1844), .Y(n4328) );
  INVX1 U3732 ( .A(n1424), .Y(n4320) );
  INVX1 U3733 ( .A(fpuReady), .Y(n4113) );
  INVX1 U3734 ( .A(n4333), .Y(n4336) );
  INVX1 U3735 ( .A(n4107), .Y(n3718) );
  OR2X1 U3736 ( .A(n2309), .B(n3549), .Y(n4110) );
  INVX1 U3737 ( .A(n3725), .Y(n4120) );
  AND2X1 U3738 ( .A(n4142), .B(n4135), .Y(n524) );
  INVX1 U3739 ( .A(n1275), .Y(n1020) );
  INVX1 U3740 ( .A(pc[17]), .Y(n1119) );
  INVX1 U3741 ( .A(pc[19]), .Y(n1117) );
  INVX1 U3742 ( .A(pc[18]), .Y(n1118) );
  INVX1 U3743 ( .A(pc[20]), .Y(n1116) );
  INVX1 U3744 ( .A(pc[16]), .Y(n1120) );
  INVX1 U3745 ( .A(pc[24]), .Y(n1112) );
  INVX1 U3746 ( .A(pc[21]), .Y(n1115) );
  INVX1 U3747 ( .A(pc[22]), .Y(n1114) );
  INVX1 U3748 ( .A(pc[26]), .Y(n1110) );
  INVX1 U3749 ( .A(pc[23]), .Y(n1113) );
  INVX1 U3750 ( .A(pc[27]), .Y(n1109) );
  INVX1 U3751 ( .A(pc[28]), .Y(n1108) );
  INVX1 U3752 ( .A(pc[25]), .Y(n1111) );
  INVX1 U3753 ( .A(pc[29]), .Y(n1107) );
  INVX1 U3754 ( .A(pc[30]), .Y(n1106) );
  INVX1 U3755 ( .A(pc[31]), .Y(n1105) );
  INVX1 U3756 ( .A(pc[6]), .Y(n4348) );
  INVX1 U3757 ( .A(pc[7]), .Y(n4349) );
  INVX1 U3758 ( .A(pc[9]), .Y(n4351) );
  INVX1 U3759 ( .A(pc[8]), .Y(n4350) );
  INVX1 U3760 ( .A(pc[14]), .Y(n4356) );
  INVX1 U3761 ( .A(pc[3]), .Y(n4345) );
  INVX1 U3762 ( .A(pc[13]), .Y(n4355) );
  INVX1 U3763 ( .A(pc[4]), .Y(n4346) );
  INVX1 U3764 ( .A(pc[12]), .Y(n4354) );
  INVX1 U3765 ( .A(pc[10]), .Y(n4352) );
  INVX1 U3766 ( .A(pc[1]), .Y(n4343) );
  INVX1 U3767 ( .A(pc[15]), .Y(n4357) );
  INVX1 U3768 ( .A(pc[2]), .Y(n4344) );
  INVX1 U3769 ( .A(pc[0]), .Y(n4342) );
  INVX1 U3770 ( .A(pc[5]), .Y(n4347) );
  INVX1 U3771 ( .A(pc[11]), .Y(n4353) );
  INVX1 U3772 ( .A(N1161), .Y(n589) );
  INVX1 U3773 ( .A(N1162), .Y(n590) );
  INVX1 U3774 ( .A(N1164), .Y(n591) );
  INVX1 U3775 ( .A(N1165), .Y(n592) );
  INVX1 U3776 ( .A(N1176), .Y(n599) );
  INVX1 U3777 ( .A(N1137), .Y(n573) );
  INVX1 U3778 ( .A(N1177), .Y(n600) );
  INVX1 U3779 ( .A(N1138), .Y(n574) );
  OR2X1 U3780 ( .A(n4174), .B(n4173), .Y(n855) );
  INVX1 U3781 ( .A(N1182), .Y(n603) );
  INVX1 U3782 ( .A(N1143), .Y(n577) );
  INVX1 U3783 ( .A(N1179), .Y(n601) );
  INVX1 U3784 ( .A(N1188), .Y(n607) );
  INVX1 U3785 ( .A(N1140), .Y(n575) );
  INVX1 U3786 ( .A(N1185), .Y(n605) );
  INVX1 U3787 ( .A(N1186), .Y(n606) );
  INVX1 U3788 ( .A(n3564), .Y(n1461) );
  INVX1 U3789 ( .A(N1183), .Y(n604) );
  INVX1 U3790 ( .A(N1147), .Y(n580) );
  INVX1 U3791 ( .A(N1146), .Y(n579) );
  OR2X1 U3792 ( .A(n4170), .B(n4173), .Y(n849) );
  INVX1 U3793 ( .A(N1149), .Y(n581) );
  INVX1 U3794 ( .A(n4315), .Y(n1462) );
  INVX1 U3795 ( .A(N1144), .Y(n578) );
  OR2X1 U3796 ( .A(n4171), .B(n4173), .Y(n851) );
  INVX1 U3797 ( .A(N1180), .Y(n602) );
  INVX1 U3798 ( .A(N1189), .Y(n608) );
  INVX1 U3799 ( .A(n4294), .Y(n1460) );
  INVX1 U3800 ( .A(n4304), .Y(n1459) );
  INVX1 U3801 ( .A(N1141), .Y(n576) );
  OR2X1 U3802 ( .A(n4172), .B(n4173), .Y(n853) );
  INVX1 U3803 ( .A(n4316), .Y(n1463) );
  INVX1 U3804 ( .A(n3563), .Y(n1464) );
  INVX1 U3805 ( .A(N1150), .Y(n582) );
  INVX1 U3806 ( .A(n4308), .Y(n1481) );
  INVX1 U3807 ( .A(n4296), .Y(n1469) );
  INVX1 U3808 ( .A(n4297), .Y(n1470) );
  INVX1 U3809 ( .A(n4309), .Y(n1482) );
  INVX1 U3810 ( .A(n4341), .Y(n1458) );
  INVX1 U3811 ( .A(n4299), .Y(n1472) );
  INVX1 U3812 ( .A(n4300), .Y(n1473) );
  INVX1 U3813 ( .A(n4318), .Y(n1465) );
  INVX1 U3814 ( .A(n4307), .Y(n1480) );
  INVX1 U3815 ( .A(n4306), .Y(n1479) );
  INVX1 U3816 ( .A(n4310), .Y(n1483) );
  INVX1 U3817 ( .A(n4301), .Y(n1475) );
  INVX1 U3818 ( .A(n4295), .Y(n1468) );
  INVX1 U3819 ( .A(n4298), .Y(n1471) );
  INVX1 U3820 ( .A(n4305), .Y(n1478) );
  INVX1 U3821 ( .A(n4181), .Y(n4177) );
  INVX1 U3822 ( .A(ir[20]), .Y(n4175) );
  INVX1 U3823 ( .A(n4319), .Y(n1467) );
  INVX1 U3824 ( .A(n4303), .Y(n1477) );
  INVX1 U3825 ( .A(n4302), .Y(n1476) );
  INVX1 U3826 ( .A(N1129), .Y(n568) );
  INVX1 U3827 ( .A(N1126), .Y(n566) );
  INVX1 U3828 ( .A(n4311), .Y(n1484) );
  INVX1 U3829 ( .A(N1128), .Y(n567) );
  INVX1 U3830 ( .A(N1125), .Y(n565) );
  INVX1 U3831 ( .A(N1135), .Y(n572) );
  INVX1 U3832 ( .A(N1132), .Y(n570) );
  INVX1 U3833 ( .A(n4159), .Y(n4160) );
  INVX1 U3834 ( .A(N1134), .Y(n571) );
  INVX1 U3835 ( .A(N1123), .Y(n564) );
  INVX1 U3836 ( .A(n4312), .Y(n1485) );
  INVX1 U3837 ( .A(N1117), .Y(n560) );
  INVX1 U3838 ( .A(N1131), .Y(n569) );
  INVX1 U3839 ( .A(N1122), .Y(n563) );
  INVX1 U3840 ( .A(N1116), .Y(n559) );
  INVX1 U3841 ( .A(n4158), .Y(n553) );
  INVX1 U3842 ( .A(aluOperand1[24]), .Y(n4257) );
  INVX1 U3843 ( .A(n4161), .Y(n4148) );
  INVX1 U3844 ( .A(N1120), .Y(n562) );
  INVX1 U3845 ( .A(aluOperand1[22]), .Y(n4242) );
  INVX1 U3846 ( .A(N1119), .Y(n561) );
  INVX1 U3847 ( .A(aluOperand1[21]), .Y(n4234) );
  INVX1 U3848 ( .A(N1206), .Y(n619) );
  INVX1 U3849 ( .A(n3281), .Y(n4021) );
  INVX1 U3850 ( .A(N1209), .Y(n621) );
  INVX1 U3851 ( .A(n3738), .Y(n3766) );
  INVX1 U3852 ( .A(n3168), .Y(n3767) );
  INVX1 U3853 ( .A(N1210), .Y(n622) );
  INVX1 U3854 ( .A(N1207), .Y(n620) );
  INVX1 U3855 ( .A(n3272), .Y(n3901) );
  INVX1 U3856 ( .A(n3269), .Y(n3904) );
  INVX1 U3857 ( .A(n3279), .Y(n4020) );
  INVX1 U3858 ( .A(N1170), .Y(n595) );
  INVX1 U3859 ( .A(n4313), .Y(n1487) );
  INVX1 U3860 ( .A(N1167), .Y(n593) );
  INVX1 U3861 ( .A(n3274), .Y(n4016) );
  INVX1 U3862 ( .A(n3271), .Y(n3905) );
  INVX1 U3863 ( .A(n3270), .Y(n3900) );
  INVX1 U3864 ( .A(n3964), .Y(\arithmetic_logic_unit/N284 ) );
  INVX1 U3865 ( .A(N1171), .Y(n596) );
  INVX1 U3866 ( .A(n3268), .Y(n3902) );
  INVX1 U3867 ( .A(N1168), .Y(n594) );
  INVX1 U3868 ( .A(N1173), .Y(n597) );
  INVX1 U3869 ( .A(n3276), .Y(n4019) );
  INVX1 U3870 ( .A(n3924), .Y(n4018) );
  INVX1 U3871 ( .A(n1843), .Y(n4155) );
  INVX1 U3872 ( .A(n3560), .Y(n4163) );
  OR2X1 U3873 ( .A(n3549), .B(n3719), .Y(n4153) );
  INVX1 U3874 ( .A(n3275), .Y(n4017) );
  INVX1 U3875 ( .A(n3915), .Y(n4015) );
  INVX1 U3876 ( .A(n3273), .Y(n3903) );
  INVX1 U3877 ( .A(N1203), .Y(n617) );
  INVX1 U3878 ( .A(N1174), .Y(n598) );
  INVX1 U3879 ( .A(N1197), .Y(n613) );
  INVX1 U3880 ( .A(N1191), .Y(n609) );
  INVX1 U3881 ( .A(N1201), .Y(n616) );
  INVX1 U3882 ( .A(N1192), .Y(n610) );
  INVX1 U3883 ( .A(N1204), .Y(n618) );
  AND2X1 U3884 ( .A(n4130), .B(n3724), .Y(n4333) );
  INVX1 U3885 ( .A(n4130), .Y(n4136) );
  INVX1 U3886 ( .A(n2404), .Y(n4107) );
  INVX1 U3887 ( .A(opcode[2]), .Y(n4329) );
  INVX1 U3888 ( .A(n2413), .Y(n4115) );
  INVX1 U3889 ( .A(opcode[5]), .Y(n4105) );
  INVX1 U3890 ( .A(n1849), .Y(n4145) );
  INVX1 U3891 ( .A(aluOperation[2]), .Y(n4369) );
  INVX1 U3892 ( .A(n3685), .Y(n3911) );
  AND2X1 U3893 ( .A(n4368), .B(aluOperation[2]), .Y(n4104) );
  INVX1 U3894 ( .A(aluOperation[1]), .Y(n4368) );
  INVX1 U3895 ( .A(n3240), .Y(\lt_x_1100_4/B[26] ) );
  INVX1 U3896 ( .A(aluSrcB[1]), .Y(n4100) );
  INVX1 U3897 ( .A(aluSrcA[0]), .Y(n4035) );
  INVX1 U3898 ( .A(aluSrcB[0]), .Y(n4092) );
  INVX1 U3899 ( .A(reset), .Y(n4364) );
  INVX1 U3900 ( .A(n3670), .Y(\sub_x_1100_2/B[4] ) );
  BUFX2 U3901 ( .A(aluOperand1[29]), .Y(\sub_x_1100_2/A[29] ) );
  BUFX2 U3902 ( .A(aluOperand1[31]), .Y(\sub_x_1100_2/A[31] ) );
  BUFX2 U3903 ( .A(aluOperand1[3]), .Y(n3721) );
  BUFX2 U3904 ( .A(aluOperand1[1]), .Y(n3722) );
  INVX1 U3905 ( .A(n3517), .Y(n4151) );
  BUFX2 U3906 ( .A(aluOperand1[30]), .Y(\sub_x_1100_2/A[30] ) );
  AND2X1 U3907 ( .A(aluOperation[3]), .B(n245), .Y(n3708) );
  BUFX2 U3908 ( .A(aluOperand1[28]), .Y(\sub_x_1100_2/A[28] ) );
  INVX1 U3909 ( .A(aluOperand1[18]), .Y(n3760) );
  INVX1 U3910 ( .A(n3650), .Y(\lt_x_1100_4/B[29] ) );
  INVX1 U3911 ( .A(\sub_x_1100_2/A[2] ), .Y(n3752) );
  INVX1 U3912 ( .A(n3283), .Y(\lt_x_1100_4/B[30] ) );
  INVX1 U3913 ( .A(n3257), .Y(\lt_x_1100_4/B[28] ) );
  INVX1 U3914 ( .A(n3282), .Y(\lt_x_1100_4/B[31] ) );
  INVX1 U3915 ( .A(n4099), .Y(\lt_x_1100_4/B[5] ) );
  INVX1 U3916 ( .A(n4097), .Y(\lt_x_1100_4/B[7] ) );
  INVX1 U3917 ( .A(n3258), .Y(\lt_x_1100_4/B[27] ) );
  INVX1 U3918 ( .A(n4213), .Y(\lt_x_1100_4/B[13] ) );
  INVX1 U3919 ( .A(n4215), .Y(\lt_x_1100_4/B[15] ) );
  INVX1 U3920 ( .A(n3248), .Y(\lt_x_1100_4/B[17] ) );
  INVX1 U3921 ( .A(n3247), .Y(\lt_x_1100_4/B[19] ) );
  INVX1 U3922 ( .A(n3243), .Y(\lt_x_1100_4/B[23] ) );
  INVX1 U3923 ( .A(n3241), .Y(\lt_x_1100_4/B[25] ) );
  INVX1 U3924 ( .A(\sub_x_1100_2/A[29] ), .Y(n3753) );
  INVX1 U3925 ( .A(n4098), .Y(\lt_x_1100_4/B[6] ) );
  INVX1 U3926 ( .A(n2292), .Y(n3765) );
  INVX1 U3927 ( .A(n4094), .Y(\lt_x_1100_4/B[10] ) );
  INVX1 U3928 ( .A(n4093), .Y(\lt_x_1100_4/B[16] ) );
  INVX1 U3929 ( .A(n1381), .Y(n4269) );
  INVX1 U3930 ( .A(n3244), .Y(\lt_x_1100_4/B[22] ) );
  INVX1 U3931 ( .A(n4096), .Y(\lt_x_1100_4/B[8] ) );
  INVX1 U3932 ( .A(n3242), .Y(\lt_x_1100_4/B[24] ) );
  INVX1 U3933 ( .A(n3246), .Y(\lt_x_1100_4/B[20] ) );
  INVX1 U3934 ( .A(n4095), .Y(\lt_x_1100_4/B[9] ) );
  INVX1 U3935 ( .A(n3245), .Y(\lt_x_1100_4/B[21] ) );
  BUFX2 U3936 ( .A(aluOperand1[27]), .Y(\sub_x_1100_2/A[27] ) );
  INVX1 U3937 ( .A(\sub_x_1100_2/A[27] ), .Y(n3754) );
  INVX1 U3938 ( .A(n3722), .Y(n3758) );
  INVX1 U3939 ( .A(n3721), .Y(n3750) );
  INVX1 U3940 ( .A(aluOperand1[17]), .Y(n3761) );
  INVX1 U3941 ( .A(\sub_x_1100_2/A[31] ), .Y(n3751) );
  INVX1 U3942 ( .A(aluOperand1[19]), .Y(n3759) );
  INVX1 U3943 ( .A(aluOperand1[23]), .Y(n3757) );
  INVX1 U3944 ( .A(aluOperand1[25]), .Y(n3756) );
  INVX1 U3945 ( .A(aluOperand1[26]), .Y(n3755) );
  INVX1 U3946 ( .A(aluOperand1[11]), .Y(n3764) );
  INVX1 U3947 ( .A(aluOperand1[13]), .Y(n3763) );
  INVX1 U3948 ( .A(n2060), .Y(n3762) );
  INVX1 U3949 ( .A(aluOperand1[5]), .Y(n3749) );
  INVX1 U3950 ( .A(aluOperand1[7]), .Y(n3748) );
  OR2X1 U3951 ( .A(pcWrite), .B(reset), .Y(n3715) );
  INVX1 U3952 ( .A(\funct3[0] ), .Y(n1145) );
  INVX1 U3953 ( .A(aluResultRegister[0]), .Y(n4090) );
  INVX1 U3954 ( .A(aluResultRegister[1]), .Y(n4088) );
  INVX1 U3955 ( .A(aluResultRegister[2]), .Y(n4086) );
  INVX1 U3956 ( .A(aluResultRegister[3]), .Y(n4084) );
  INVX1 U3957 ( .A(aluResultRegister[4]), .Y(n4082) );
  INVX1 U3958 ( .A(aluResultRegister[5]), .Y(n4080) );
  INVX1 U3959 ( .A(aluResultRegister[6]), .Y(n4078) );
  INVX1 U3960 ( .A(aluResultRegister[7]), .Y(n4076) );
  INVX1 U3961 ( .A(aluResultRegister[8]), .Y(n4074) );
  INVX1 U3962 ( .A(aluResultRegister[9]), .Y(n4072) );
  INVX1 U3963 ( .A(aluResultRegister[10]), .Y(n4070) );
  INVX1 U3964 ( .A(aluResultRegister[11]), .Y(n4068) );
  INVX1 U3965 ( .A(aluResultRegister[12]), .Y(n4066) );
  INVX1 U3966 ( .A(aluResultRegister[13]), .Y(n4064) );
  INVX1 U3967 ( .A(aluResultRegister[14]), .Y(n4062) );
  INVX1 U3968 ( .A(aluResultRegister[15]), .Y(n4060) );
  INVX1 U3969 ( .A(aluResultRegister[16]), .Y(n4058) );
  INVX1 U3970 ( .A(aluResultRegister[17]), .Y(n4056) );
  INVX1 U3971 ( .A(aluResultRegister[18]), .Y(n4054) );
  INVX1 U3972 ( .A(aluResultRegister[19]), .Y(n4052) );
  INVX1 U3973 ( .A(aluResultRegister[20]), .Y(n4050) );
  INVX1 U3974 ( .A(aluResultRegister[21]), .Y(n4048) );
  INVX1 U3975 ( .A(aluResultRegister[22]), .Y(n4046) );
  INVX1 U3976 ( .A(aluResultRegister[23]), .Y(n4044) );
  INVX1 U3977 ( .A(aluResultRegister[24]), .Y(n4042) );
  INVX1 U3978 ( .A(aluResultRegister[25]), .Y(n4040) );
  INVX1 U3979 ( .A(aluResultRegister[26]), .Y(n4038) );
  OR2X1 U3980 ( .A(reset), .B(irWrite), .Y(n3716) );
  INVX1 U3981 ( .A(funct3[2]), .Y(n4117) );
  BUFX2 U3982 ( .A(n4165), .Y(n3719) );
  INVX1 U3983 ( .A(n2290), .Y(n4326) );
  INVX1 U3984 ( .A(N1195), .Y(n612) );
  INVX1 U3985 ( .A(N1194), .Y(n611) );
  INVX1 U3986 ( .A(N1198), .Y(n614) );
  AOI22X1 U3987 ( .A(\lt_x_1100_4/B[31] ), .B(n3751), .C(\sub_x_1100_2/A[30] ), 
        .D(n3283), .Y(n3745) );
  AOI21X1 U3988 ( .A(\sub_x_1100_2/A[28] ), .B(n3257), .C(n2816), .Y(n3747) );
  AOI22X1 U3989 ( .A(n2916), .B(n2236), .C(n1831), .D(n3749), .Y(n3729) );
  AOI22X1 U3990 ( .A(\sub_x_1100_2/A[4] ), .B(n2239), .C(n1819), .D(n1858), 
        .Y(n3728) );
  AOI22X1 U3991 ( .A(n1818), .B(n2889), .C(n2286), .D(n3750), .Y(n3727) );
  AOI22X1 U3992 ( .A(n2060), .B(n1827), .C(\sub_x_1100_2/A[14] ), .D(n3250), 
        .Y(n3731) );
  AOI21X1 U3993 ( .A(\sub_x_1100_2/A[8] ), .B(n2259), .C(n3311), .Y(n3730) );
  AOI22X1 U3994 ( .A(n1846), .B(n2890), .C(\lt_x_1100_4/B[13] ), .D(n3763), 
        .Y(n3733) );
  AOI22X1 U3995 ( .A(n3249), .B(n2891), .C(\lt_x_1100_4/B[15] ), .D(n3762), 
        .Y(n3732) );
  OAI21X1 U3996 ( .A(n2875), .B(n3767), .C(n2651), .Y(n3735) );
  AOI22X1 U3997 ( .A(\lt_x_1100_4/B[10] ), .B(n2892), .C(\lt_x_1100_4/B[11] ), 
        .D(n3764), .Y(n3734) );
  AOI21X1 U3998 ( .A(aluOperand1[20]), .B(n3246), .C(n2818), .Y(n3741) );
  OAI21X1 U3999 ( .A(\lt_x_1100_4/B[18] ), .B(n3760), .C(n2254), .Y(n3738) );
  AOI22X1 U4000 ( .A(\lt_x_1100_4/B[22] ), .B(n2896), .C(\lt_x_1100_4/B[23] ), 
        .D(n3757), .Y(n3742) );
  OAI21X1 U4001 ( .A(aluOperand1[21]), .B(n3245), .C(n2227), .Y(n3736) );
  AOI22X1 U4002 ( .A(\lt_x_1100_4/B[16] ), .B(n2893), .C(\lt_x_1100_4/B[17] ), 
        .D(n3761), .Y(n3739) );
  AOI22X1 U4003 ( .A(\lt_x_1100_4/B[18] ), .B(n2897), .C(\lt_x_1100_4/B[19] ), 
        .D(n3759), .Y(n3737) );
  OAI21X1 U4004 ( .A(n2876), .B(n3738), .C(n2248), .Y(n3740) );
  AOI22X1 U4005 ( .A(\lt_x_1100_4/B[24] ), .B(n2898), .C(\lt_x_1100_4/B[25] ), 
        .D(n3756), .Y(n3744) );
  AOI22X1 U4006 ( .A(\lt_x_1100_4/B[26] ), .B(n2894), .C(\lt_x_1100_4/B[27] ), 
        .D(n3754), .Y(n3743) );
  AOI22X1 U4007 ( .A(\lt_x_1100_4/B[28] ), .B(n2895), .C(\lt_x_1100_4/B[29] ), 
        .D(n3753), .Y(n3746) );
  OAI21X1 U4008 ( .A(\lt_x_1100_4/B[26] ), .B(n3755), .C(n2234), .Y(n3790) );
  AOI22X1 U4009 ( .A(\sub_x_1100_2/A[31] ), .B(n3282), .C(\sub_x_1100_2/A[30] ), .D(n3283), .Y(n3792) );
  AOI21X1 U4010 ( .A(\sub_x_1100_2/A[28] ), .B(n3257), .C(n2820), .Y(n3793) );
  AOI22X1 U4011 ( .A(\sub_x_1100_2/A[7] ), .B(\sub_x_1100_2/n227 ), .C(
        \sub_x_1100_2/A[6] ), .D(n3765), .Y(n3773) );
  AOI21X1 U4012 ( .A(n1819), .B(n1858), .C(\sub_x_1100_2/A[4] ), .Y(n3768) );
  AOI21X1 U4013 ( .A(n3722), .B(n3910), .C(aluOperand1[0]), .Y(n3769) );
  AOI22X1 U4014 ( .A(n2917), .B(n4022), .C(\ashr_1100_6/SH[1] ), .D(n3758), 
        .Y(n3772) );
  OAI21X1 U4015 ( .A(n1818), .B(n3752), .C(n2229), .Y(n3771) );
  AOI21X1 U4016 ( .A(n3721), .B(n3712), .C(\sub_x_1100_2/A[2] ), .Y(n3770) );
  AOI21X1 U4017 ( .A(\sub_x_1100_2/A[7] ), .B(\sub_x_1100_2/n227 ), .C(
        \sub_x_1100_2/A[6] ), .Y(n3774) );
  AOI22X1 U4018 ( .A(n2293), .B(n3748), .C(n2989), .D(n2292), .Y(n3776) );
  AOI22X1 U4019 ( .A(\sub_x_1100_2/A[12] ), .B(n1856), .C(n1820), .D(n2264), 
        .Y(n3775) );
  AOI22X1 U4020 ( .A(\sub_x_1100_2/A[11] ), .B(n3252), .C(\sub_x_1100_2/A[10] ), .D(n2233), .Y(n3782) );
  AOI21X1 U4021 ( .A(n1820), .B(n2264), .C(\sub_x_1100_2/A[12] ), .Y(n3777) );
  AOI21X1 U4022 ( .A(n2060), .B(n1827), .C(\sub_x_1100_2/A[14] ), .Y(n3778) );
  AOI21X1 U4023 ( .A(\sub_x_1100_2/A[11] ), .B(n3252), .C(\sub_x_1100_2/A[10] ), .Y(n3779) );
  AOI21X1 U4024 ( .A(n2469), .B(n2260), .C(\sub_x_1100_2/A[8] ), .Y(n3780) );
  OAI21X1 U4025 ( .A(n2470), .B(n2260), .C(n2228), .Y(n3781) );
  AOI22X1 U4026 ( .A(aluOperand1[23]), .B(n3243), .C(aluOperand1[22]), .D(
        n3244), .Y(n3785) );
  AOI21X1 U4027 ( .A(aluOperand1[23]), .B(n3243), .C(aluOperand1[22]), .Y(
        n3783) );
  AOI21X1 U4028 ( .A(aluOperand1[21]), .B(n3245), .C(aluOperand1[20]), .Y(
        n3784) );
  AOI21X1 U4029 ( .A(aluOperand1[17]), .B(n2257), .C(aluOperand1[16]), .Y(
        n3786) );
  AOI21X1 U4030 ( .A(aluOperand1[19]), .B(n3247), .C(aluOperand1[18]), .Y(
        n3787) );
  AOI21X1 U4031 ( .A(aluOperand1[25]), .B(n3241), .C(aluOperand1[24]), .Y(
        n3788) );
  AOI21X1 U4032 ( .A(\sub_x_1100_2/A[27] ), .B(n3258), .C(aluOperand1[26]), 
        .Y(n3789) );
  OAI21X1 U4033 ( .A(n2244), .B(n3790), .C(n2245), .Y(n3794) );
  AOI21X1 U4034 ( .A(\sub_x_1100_2/A[29] ), .B(n3650), .C(\sub_x_1100_2/A[28] ), .Y(n3791) );
  NAND3X1 U4035 ( .A(\sub_x_1100_2/A[0] ), .B(n3910), .C(n2230), .Y(n3797) );
  AOI22X1 U4036 ( .A(n4022), .B(n3722), .C(\sub_x_1100_2/A[2] ), .D(n2193), 
        .Y(n3796) );
  AOI22X1 U4037 ( .A(n1841), .B(n2900), .C(n3381), .D(n3910), .Y(n3808) );
  AND2X1 U4038 ( .A(n2251), .B(n3354), .Y(n3824) );
  AOI22X1 U4039 ( .A(n4022), .B(n3721), .C(\sub_x_1100_2/A[4] ), .D(n3685), 
        .Y(n3795) );
  AOI22X1 U4040 ( .A(n4022), .B(\sub_x_1100_2/A[5] ), .C(\sub_x_1100_2/A[6] ), 
        .D(n2193), .Y(n3799) );
  AOI22X1 U4041 ( .A(n1841), .B(n3382), .C(n3383), .D(n3910), .Y(n3807) );
  AOI22X1 U4042 ( .A(n4022), .B(\sub_x_1100_2/A[7] ), .C(\sub_x_1100_2/A[8] ), 
        .D(n3685), .Y(n3798) );
  AOI22X1 U4043 ( .A(n4022), .B(n2470), .C(\sub_x_1100_2/A[10] ), .D(n2193), 
        .Y(n3800) );
  AOI22X1 U4044 ( .A(n1841), .B(n3385), .C(n3386), .D(n3910), .Y(n3810) );
  AOI22X1 U4045 ( .A(n2238), .B(n3384), .C(n3387), .D(n2251), .Y(n3827) );
  AOI22X1 U4046 ( .A(n2286), .B(n3824), .C(n3902), .D(n3908), .Y(n3869) );
  AOI22X1 U4047 ( .A(n4022), .B(aluOperand1[0]), .C(n3722), .D(n3685), .Y(
        n3801) );
  AOI22X1 U4048 ( .A(n4022), .B(\sub_x_1100_2/A[2] ), .C(n3721), .D(n3685), 
        .Y(n3803) );
  AOI22X1 U4049 ( .A(\ashr_1100_6/SH[1] ), .B(n3363), .C(n3388), .D(n3910), 
        .Y(n3812) );
  AND2X1 U4050 ( .A(n2251), .B(n3355), .Y(n3828) );
  AOI22X1 U4051 ( .A(n4022), .B(\sub_x_1100_2/A[4] ), .C(n1819), .D(n2193), 
        .Y(n3802) );
  AOI22X1 U4052 ( .A(n4022), .B(\sub_x_1100_2/A[6] ), .C(\sub_x_1100_2/A[7] ), 
        .D(n2193), .Y(n3805) );
  AOI22X1 U4053 ( .A(\ashr_1100_6/SH[1] ), .B(n3389), .C(n3390), .D(n3910), 
        .Y(n3811) );
  AOI22X1 U4054 ( .A(n4022), .B(\sub_x_1100_2/A[8] ), .C(n2469), .D(n2193), 
        .Y(n3804) );
  AOI22X1 U4055 ( .A(n4022), .B(\sub_x_1100_2/A[10] ), .C(\sub_x_1100_2/A[11] ), .D(n2193), .Y(n3806) );
  AOI22X1 U4056 ( .A(n1841), .B(n3392), .C(n3393), .D(n3910), .Y(n3814) );
  AOI22X1 U4057 ( .A(n2238), .B(n3391), .C(n3394), .D(n2251), .Y(n3831) );
  AOI22X1 U4058 ( .A(n3909), .B(n3828), .C(n3904), .D(n3908), .Y(n3875) );
  AOI22X1 U4059 ( .A(n1841), .B(n3381), .C(n3382), .D(n3910), .Y(n3816) );
  AOI22X1 U4060 ( .A(n2238), .B(n3364), .C(n3900), .D(n2251), .Y(n3832) );
  AOI22X1 U4061 ( .A(n1841), .B(n3383), .C(n3385), .D(n3910), .Y(n3815) );
  AOI22X1 U4062 ( .A(n2226), .B(\sub_x_1100_2/A[11] ), .C(\sub_x_1100_2/A[12] ), .D(n2230), .Y(n3809) );
  AOI22X1 U4063 ( .A(n1841), .B(n3386), .C(n3396), .D(n3910), .Y(n3818) );
  AOI22X1 U4064 ( .A(n2238), .B(n3395), .C(n3397), .D(n3906), .Y(n3835) );
  AOI22X1 U4065 ( .A(n3909), .B(n3299), .C(n3905), .D(n3908), .Y(n3882) );
  AOI22X1 U4066 ( .A(n1841), .B(n3388), .C(n3389), .D(n3910), .Y(n3820) );
  AOI22X1 U4067 ( .A(n2238), .B(n3323), .C(n3398), .D(n2251), .Y(n3836) );
  AOI22X1 U4068 ( .A(n1841), .B(n3390), .C(n3392), .D(n3910), .Y(n3819) );
  AOI22X1 U4069 ( .A(n4022), .B(\sub_x_1100_2/A[12] ), .C(n1820), .D(n2230), 
        .Y(n3813) );
  AOI22X1 U4070 ( .A(n1841), .B(n3393), .C(n3400), .D(n3910), .Y(n3822) );
  AOI22X1 U4071 ( .A(n2238), .B(n3399), .C(n3401), .D(n3906), .Y(n3839) );
  AOI22X1 U4072 ( .A(n3909), .B(n3370), .C(n3402), .D(n3908), .Y(n3886) );
  AOI22X1 U4073 ( .A(n2238), .B(n3354), .C(n3384), .D(n2251), .Y(n3841) );
  AOI22X1 U4074 ( .A(n2226), .B(n1820), .C(\sub_x_1100_2/A[14] ), .D(n2193), 
        .Y(n3817) );
  AOI22X1 U4075 ( .A(n1841), .B(n3396), .C(n3403), .D(n3910), .Y(n3826) );
  AOI22X1 U4076 ( .A(n2238), .B(n3387), .C(n3404), .D(n2251), .Y(n3844) );
  AOI22X1 U4077 ( .A(n3909), .B(n3371), .C(n3405), .D(n3908), .Y(n3890) );
  AOI22X1 U4078 ( .A(n2238), .B(n3355), .C(n3391), .D(n3906), .Y(n3846) );
  AOI22X1 U4079 ( .A(n4022), .B(\sub_x_1100_2/A[14] ), .C(n2060), .D(n2193), 
        .Y(n3821) );
  AOI22X1 U4080 ( .A(n1841), .B(n3400), .C(n3406), .D(n3910), .Y(n3830) );
  AOI22X1 U4081 ( .A(n2238), .B(n3394), .C(n3407), .D(n3906), .Y(n3849) );
  AOI22X1 U4082 ( .A(n3909), .B(n3372), .C(n3408), .D(n3908), .Y(n3894) );
  AND2X1 U4083 ( .A(n2239), .B(n3358), .Y(\arithmetic_logic_unit/N266 ) );
  AOI22X1 U4084 ( .A(n2238), .B(n3270), .C(n3395), .D(n2251), .Y(n3851) );
  AOI22X1 U4085 ( .A(n2226), .B(n2060), .C(aluOperand1[16]), .D(n2230), .Y(
        n3825) );
  AOI22X1 U4086 ( .A(n1841), .B(n3403), .C(n3409), .D(n3910), .Y(n3834) );
  AOI22X1 U4087 ( .A(n2238), .B(n3397), .C(n3410), .D(n2251), .Y(n3855) );
  AND2X1 U4088 ( .A(n3323), .B(n3906), .Y(n3858) );
  AOI22X1 U4089 ( .A(n2238), .B(n3398), .C(n3399), .D(n2251), .Y(n3857) );
  AOI22X1 U4090 ( .A(n4022), .B(aluOperand1[16]), .C(aluOperand1[17]), .D(
        n2230), .Y(n3829) );
  AOI22X1 U4091 ( .A(n1841), .B(n3406), .C(n3412), .D(n3910), .Y(n3838) );
  AOI22X1 U4092 ( .A(n2238), .B(n3401), .C(n3413), .D(n3906), .Y(n3862) );
  AOI22X1 U4093 ( .A(n3909), .B(n3273), .C(n3414), .D(n3908), .Y(n3823) );
  OAI21X1 U4094 ( .A(n3340), .B(n2239), .C(n2692), .Y(
        \arithmetic_logic_unit/N268 ) );
  AOI22X1 U4095 ( .A(n2226), .B(aluOperand1[17]), .C(aluOperand1[18]), .D(
        n2230), .Y(n3833) );
  AOI22X1 U4096 ( .A(n1841), .B(n3409), .C(n3415), .D(n3910), .Y(n3843) );
  AOI22X1 U4097 ( .A(n2238), .B(n3404), .C(n3416), .D(n2251), .Y(n3867) );
  AOI22X1 U4098 ( .A(n4022), .B(aluOperand1[18]), .C(aluOperand1[19]), .D(
        n2230), .Y(n3837) );
  AOI22X1 U4099 ( .A(n1841), .B(n3412), .C(n3418), .D(n3910), .Y(n3848) );
  AOI22X1 U4100 ( .A(n2238), .B(n3407), .C(n3419), .D(n2251), .Y(n3873) );
  AOI22X1 U4101 ( .A(n4022), .B(aluOperand1[19]), .C(aluOperand1[20]), .D(
        n2230), .Y(n3842) );
  AOI22X1 U4102 ( .A(n1841), .B(n3415), .C(n3421), .D(n3910), .Y(n3853) );
  AOI22X1 U4103 ( .A(n2238), .B(n3410), .C(n3422), .D(n3906), .Y(n3880) );
  OR2X1 U4104 ( .A(n3909), .B(n3370), .Y(n3895) );
  AOI22X1 U4105 ( .A(n3911), .B(aluOperand1[20]), .C(aluOperand1[21]), .D(
        n2230), .Y(n3847) );
  AOI22X1 U4106 ( .A(n1841), .B(n3418), .C(n3424), .D(n3910), .Y(n3860) );
  AOI22X1 U4107 ( .A(n2238), .B(n3413), .C(n3425), .D(n3906), .Y(n3885) );
  AOI22X1 U4108 ( .A(n3909), .B(n3402), .C(n3426), .D(n3908), .Y(n3840) );
  OAI21X1 U4109 ( .A(n3895), .B(n2239), .C(n2693), .Y(
        \arithmetic_logic_unit/N272 ) );
  OR2X1 U4110 ( .A(n3909), .B(n3371), .Y(n3896) );
  AOI22X1 U4111 ( .A(n4022), .B(aluOperand1[21]), .C(aluOperand1[22]), .D(
        n2230), .Y(n3852) );
  AOI22X1 U4112 ( .A(n1841), .B(n3421), .C(n3427), .D(n3910), .Y(n3865) );
  AOI22X1 U4113 ( .A(n2238), .B(n3416), .C(n3428), .D(n3906), .Y(n3889) );
  AOI22X1 U4114 ( .A(n3909), .B(n3405), .C(n3429), .D(n3908), .Y(n3845) );
  OAI21X1 U4115 ( .A(n3896), .B(n2239), .C(n2694), .Y(
        \arithmetic_logic_unit/N273 ) );
  OR2X1 U4116 ( .A(n3909), .B(n3372), .Y(n3897) );
  AOI22X1 U4117 ( .A(n4022), .B(aluOperand1[22]), .C(aluOperand1[23]), .D(
        n2193), .Y(n3859) );
  AOI22X1 U4118 ( .A(n1841), .B(n3424), .C(n3430), .D(n3910), .Y(n3871) );
  AOI22X1 U4119 ( .A(n2238), .B(n3419), .C(n3431), .D(n3906), .Y(n3893) );
  AOI22X1 U4120 ( .A(n3909), .B(n3408), .C(n3432), .D(n3908), .Y(n3850) );
  OAI21X1 U4121 ( .A(n3897), .B(n2239), .C(n2385), .Y(
        \arithmetic_logic_unit/N274 ) );
  AOI22X1 U4122 ( .A(n3909), .B(n3290), .C(n3901), .D(n3908), .Y(n3898) );
  AOI22X1 U4123 ( .A(n3911), .B(aluOperand1[23]), .C(aluOperand1[24]), .D(
        n2230), .Y(n3864) );
  AOI22X1 U4124 ( .A(n1841), .B(n3427), .C(n3433), .D(n3910), .Y(n3878) );
  AOI22X1 U4125 ( .A(n2238), .B(n3422), .C(n3434), .D(n3906), .Y(n3854) );
  AOI22X1 U4126 ( .A(n3909), .B(n3411), .C(n2974), .D(n3908), .Y(n3856) );
  OAI21X1 U4127 ( .A(n3329), .B(n2239), .C(n2695), .Y(
        \arithmetic_logic_unit/N275 ) );
  AOI22X1 U4128 ( .A(n3909), .B(n3858), .C(n3903), .D(n3908), .Y(n3899) );
  AOI22X1 U4129 ( .A(n3911), .B(aluOperand1[24]), .C(aluOperand1[25]), .D(
        n2230), .Y(n3870) );
  AOI22X1 U4130 ( .A(n1841), .B(n3430), .C(n3435), .D(n3910), .Y(n3884) );
  AOI22X1 U4131 ( .A(n2238), .B(n3425), .C(n3436), .D(n3906), .Y(n3861) );
  AOI22X1 U4132 ( .A(n3909), .B(n3414), .C(n2975), .D(n3908), .Y(n3863) );
  OAI21X1 U4133 ( .A(n3330), .B(n2239), .C(n2696), .Y(
        \arithmetic_logic_unit/N276 ) );
  AOI22X1 U4134 ( .A(n4022), .B(aluOperand1[25]), .C(aluOperand1[26]), .D(
        n2230), .Y(n3876) );
  AOI22X1 U4135 ( .A(n1841), .B(n3433), .C(n3437), .D(n3910), .Y(n3888) );
  AOI22X1 U4136 ( .A(n2238), .B(n3428), .C(n3438), .D(n3906), .Y(n3866) );
  AOI22X1 U4137 ( .A(n3909), .B(n3417), .C(n2976), .D(n3908), .Y(n3868) );
  OAI21X1 U4138 ( .A(n3326), .B(n2239), .C(n2697), .Y(
        \arithmetic_logic_unit/N277 ) );
  AOI22X1 U4139 ( .A(n4022), .B(aluOperand1[26]), .C(\sub_x_1100_2/A[27] ), 
        .D(n2230), .Y(n3883) );
  AOI22X1 U4140 ( .A(n1841), .B(n3435), .C(n3439), .D(n3910), .Y(n3892) );
  AOI22X1 U4141 ( .A(n2238), .B(n3431), .C(n3440), .D(n3906), .Y(n3872) );
  AOI22X1 U4142 ( .A(n3909), .B(n3420), .C(n2977), .D(n3908), .Y(n3874) );
  OAI21X1 U4143 ( .A(n3327), .B(n2239), .C(n2699), .Y(
        \arithmetic_logic_unit/N278 ) );
  AOI22X1 U4144 ( .A(n4022), .B(\sub_x_1100_2/A[27] ), .C(\sub_x_1100_2/A[28] ), .D(n2230), .Y(n3887) );
  AOI22X1 U4145 ( .A(n1841), .B(n3437), .C(n3441), .D(n3910), .Y(n3877) );
  AOI22X1 U4146 ( .A(n2238), .B(n3434), .C(n2978), .D(n3906), .Y(n3879) );
  AOI22X1 U4147 ( .A(n3909), .B(n3423), .C(n2979), .D(n3908), .Y(n3881) );
  OAI21X1 U4148 ( .A(n3328), .B(n2239), .C(n2308), .Y(
        \arithmetic_logic_unit/N279 ) );
  AOI22X1 U4149 ( .A(n1823), .B(\sub_x_1100_2/A[28] ), .C(\sub_x_1100_2/A[29] ), .D(n2193), .Y(n3891) );
  AOI22X1 U4150 ( .A(n4022), .B(\sub_x_1100_2/A[31] ), .C(\sub_x_1100_2/A[30] ), .D(n3685), .Y(n3912) );
  AOI22X1 U4151 ( .A(n4022), .B(\sub_x_1100_2/A[29] ), .C(\sub_x_1100_2/A[28] ), .D(n2193), .Y(n3914) );
  AOI22X1 U4152 ( .A(\ashr_1100_6/SH[1] ), .B(n3373), .C(n3443), .D(n3910), 
        .Y(n3965) );
  AOI22X1 U4153 ( .A(n4022), .B(\sub_x_1100_2/A[27] ), .C(aluOperand1[26]), 
        .D(n2193), .Y(n3913) );
  AOI22X1 U4154 ( .A(n4022), .B(aluOperand1[25]), .C(aluOperand1[24]), .D(
        n2193), .Y(n3917) );
  AOI22X1 U4155 ( .A(n1841), .B(n3444), .C(n3445), .D(n3910), .Y(n3927) );
  AOI22X1 U4156 ( .A(n2238), .B(n3550), .C(n3446), .D(n2251), .Y(n3971) );
  AOI22X1 U4157 ( .A(n4022), .B(aluOperand1[23]), .C(aluOperand1[22]), .D(
        n2193), .Y(n3916) );
  AOI22X1 U4158 ( .A(n4022), .B(aluOperand1[21]), .C(aluOperand1[20]), .D(
        n2193), .Y(n3919) );
  AOI22X1 U4159 ( .A(n1841), .B(n3447), .C(n3448), .D(n3910), .Y(n3926) );
  AOI22X1 U4160 ( .A(n4022), .B(aluOperand1[19]), .C(aluOperand1[18]), .D(
        n3685), .Y(n3918) );
  AOI22X1 U4161 ( .A(n4022), .B(aluOperand1[17]), .C(aluOperand1[16]), .D(
        n3685), .Y(n3921) );
  AOI22X1 U4162 ( .A(n1841), .B(n3450), .C(n3451), .D(n3910), .Y(n3929) );
  AOI22X1 U4163 ( .A(n2238), .B(n3449), .C(n3452), .D(n2251), .Y(n4010) );
  AOI22X1 U4164 ( .A(n2286), .B(n3374), .C(n3453), .D(n3908), .Y(n3948) );
  AOI22X1 U4165 ( .A(n4022), .B(n2060), .C(\sub_x_1100_2/A[14] ), .D(n2193), 
        .Y(n3920) );
  AOI22X1 U4166 ( .A(n4022), .B(n1820), .C(\sub_x_1100_2/A[12] ), .D(n2193), 
        .Y(n3923) );
  AOI22X1 U4167 ( .A(n1841), .B(n3454), .C(n3455), .D(n3910), .Y(n3928) );
  AOI22X1 U4168 ( .A(n4022), .B(\sub_x_1100_2/A[11] ), .C(\sub_x_1100_2/A[10] ), .D(n2193), .Y(n3922) );
  AOI22X1 U4169 ( .A(n4022), .B(n2469), .C(\sub_x_1100_2/A[8] ), .D(n2193), 
        .Y(n3975) );
  AOI22X1 U4170 ( .A(n1841), .B(n3457), .C(n3458), .D(n3910), .Y(n3990) );
  AOI22X1 U4171 ( .A(n2238), .B(n3456), .C(n3459), .D(n2251), .Y(n4009) );
  AOI22X1 U4172 ( .A(n4022), .B(\sub_x_1100_2/A[7] ), .C(\sub_x_1100_2/A[6] ), 
        .D(n3685), .Y(n3974) );
  AOI22X1 U4173 ( .A(n4022), .B(n1819), .C(\sub_x_1100_2/A[4] ), .D(n2230), 
        .Y(n3977) );
  AOI22X1 U4174 ( .A(n1841), .B(n3461), .C(n3462), .D(n3910), .Y(n3989) );
  AOI22X1 U4175 ( .A(n4022), .B(n3721), .C(\sub_x_1100_2/A[2] ), .D(n3685), 
        .Y(n3976) );
  OR2X1 U4176 ( .A(n1841), .B(n3373), .Y(n3939) );
  AOI22X1 U4177 ( .A(\ashr_1100_6/SH[1] ), .B(n3443), .C(n3444), .D(n3910), 
        .Y(n3915) );
  AOI22X1 U4178 ( .A(n2238), .B(n3939), .C(n4015), .D(n2251), .Y(n3954) );
  AOI22X1 U4179 ( .A(n1841), .B(n3445), .C(n3447), .D(n3910), .Y(n3940) );
  AOI22X1 U4180 ( .A(n1841), .B(n3448), .C(n3450), .D(n3910), .Y(n3942) );
  AOI22X1 U4181 ( .A(n2238), .B(n3274), .C(n3465), .D(n2251), .Y(n3953) );
  AOI22X1 U4182 ( .A(\ashr_1100_6/SH[1] ), .B(n3451), .C(n3454), .D(n3910), 
        .Y(n3941) );
  AOI22X1 U4183 ( .A(n1841), .B(n3455), .C(n3457), .D(n3910), .Y(n4000) );
  AOI22X1 U4184 ( .A(n2238), .B(n3466), .C(n3467), .D(n2251), .Y(n3978) );
  NAND3X1 U4185 ( .A(\sub_x_1100_2/A[31] ), .B(n3910), .C(n2193), .Y(n3943) );
  AOI22X1 U4186 ( .A(n4022), .B(\sub_x_1100_2/A[30] ), .C(\sub_x_1100_2/A[29] ), .D(n2193), .Y(n3930) );
  AOI22X1 U4187 ( .A(n4022), .B(\sub_x_1100_2/A[28] ), .C(\sub_x_1100_2/A[27] ), .D(n3685), .Y(n3932) );
  AOI22X1 U4188 ( .A(n1841), .B(n3469), .C(n3470), .D(n3910), .Y(n3924) );
  AOI22X1 U4189 ( .A(n2238), .B(n3365), .C(n4018), .D(n2251), .Y(n3956) );
  AOI22X1 U4190 ( .A(n4022), .B(aluOperand1[26]), .C(aluOperand1[25]), .D(
        n2193), .Y(n3931) );
  AOI22X1 U4191 ( .A(n4022), .B(aluOperand1[24]), .C(aluOperand1[23]), .D(
        n3685), .Y(n3934) );
  AOI22X1 U4192 ( .A(n1841), .B(n3471), .C(n3472), .D(n3910), .Y(n3944) );
  AOI22X1 U4193 ( .A(n4022), .B(aluOperand1[22]), .C(aluOperand1[21]), .D(
        n3685), .Y(n3933) );
  AOI22X1 U4194 ( .A(n4022), .B(aluOperand1[20]), .C(aluOperand1[19]), .D(
        n2193), .Y(n3936) );
  AOI22X1 U4195 ( .A(\ashr_1100_6/SH[1] ), .B(n3473), .C(n3474), .D(n3910), 
        .Y(n3946) );
  AOI22X1 U4196 ( .A(n2238), .B(n3276), .C(n3475), .D(n2251), .Y(n3955) );
  AOI22X1 U4197 ( .A(n4022), .B(aluOperand1[18]), .C(aluOperand1[17]), .D(
        n2193), .Y(n3935) );
  AOI22X1 U4198 ( .A(n4022), .B(aluOperand1[16]), .C(n2060), .D(n3685), .Y(
        n3938) );
  AOI22X1 U4199 ( .A(n1841), .B(n3476), .C(n3477), .D(n3910), .Y(n3945) );
  AOI22X1 U4200 ( .A(n4022), .B(\sub_x_1100_2/A[14] ), .C(n1820), .D(n2193), 
        .Y(n3937) );
  AOI22X1 U4201 ( .A(n4022), .B(\sub_x_1100_2/A[12] ), .C(\sub_x_1100_2/A[11] ), .D(n2193), .Y(n3957) );
  AOI22X1 U4202 ( .A(n1841), .B(n3479), .C(n3480), .D(n3910), .Y(n4006) );
  AOI22X1 U4203 ( .A(n2238), .B(n3478), .C(n3481), .D(n2251), .Y(n3986) );
  AOI22X1 U4204 ( .A(n2286), .B(n3278), .C(n3482), .D(n3908), .Y(n3925) );
  OAI21X1 U4205 ( .A(n3350), .B(n2239), .C(n2701), .Y(
        \arithmetic_logic_unit/N294 ) );
  NAND3X1 U4206 ( .A(n3908), .B(n2251), .C(n3550), .Y(n3973) );
  AOI22X1 U4207 ( .A(n2238), .B(n3446), .C(n3449), .D(n2251), .Y(n3966) );
  AOI22X1 U4208 ( .A(n2238), .B(n3452), .C(n3456), .D(n2251), .Y(n3991) );
  AOI22X1 U4209 ( .A(n1841), .B(n2906), .C(n3469), .D(n3910), .Y(n3950) );
  AND2X1 U4210 ( .A(n2251), .B(n3360), .Y(n3968) );
  AOI22X1 U4211 ( .A(n1841), .B(n3470), .C(n3471), .D(n3910), .Y(n3949) );
  AOI22X1 U4212 ( .A(n1841), .B(n3472), .C(n3473), .D(n3910), .Y(n3952) );
  AOI22X1 U4213 ( .A(n2238), .B(n3485), .C(n3486), .D(n2251), .Y(n3967) );
  AOI22X1 U4214 ( .A(n1841), .B(n3474), .C(n3476), .D(n3910), .Y(n3951) );
  AOI22X1 U4215 ( .A(n1841), .B(n3477), .C(n3479), .D(n3910), .Y(n3958) );
  AOI22X1 U4216 ( .A(n2238), .B(n3487), .C(n3488), .D(n2251), .Y(n3996) );
  AOI22X1 U4217 ( .A(n2238), .B(n4015), .C(n4016), .D(n2251), .Y(n3969) );
  AOI22X1 U4218 ( .A(n2238), .B(n3465), .C(n3466), .D(n2251), .Y(n4002) );
  AOI22X1 U4219 ( .A(n2238), .B(n4018), .C(n4019), .D(n2251), .Y(n3970) );
  AOI22X1 U4220 ( .A(n2238), .B(n3475), .C(n3478), .D(n2251), .Y(n4007) );
  AOI22X1 U4221 ( .A(n2286), .B(n3491), .C(n4021), .D(n3908), .Y(n3947) );
  AOI22X1 U4222 ( .A(n2236), .B(n3368), .C(n2980), .D(n2239), .Y(
        \arithmetic_logic_unit/N298 ) );
  AOI22X1 U4223 ( .A(n2238), .B(n3360), .C(n3485), .D(n2251), .Y(n3972) );
  AOI22X1 U4224 ( .A(n2238), .B(n3486), .C(n3487), .D(n2251), .Y(n4013) );
  AOI22X1 U4225 ( .A(n2286), .B(n3375), .C(n3492), .D(n3908), .Y(n3963) );
  AND2X1 U4226 ( .A(n2239), .B(n3361), .Y(\arithmetic_logic_unit/N300 ) );
  AOI22X1 U4227 ( .A(n2286), .B(n3300), .C(n4017), .D(n3908), .Y(n3979) );
  AOI22X1 U4228 ( .A(n2286), .B(n3301), .C(n3277), .D(n3908), .Y(n3988) );
  AOI22X1 U4229 ( .A(n4022), .B(\sub_x_1100_2/A[10] ), .C(n2470), .D(n2193), 
        .Y(n3981) );
  AOI22X1 U4230 ( .A(n1841), .B(n3480), .C(n3493), .D(n3910), .Y(n3994) );
  AOI22X1 U4231 ( .A(n2238), .B(n3488), .C(n3494), .D(n2251), .Y(n4012) );
  AOI22X1 U4232 ( .A(n4022), .B(\sub_x_1100_2/A[8] ), .C(\sub_x_1100_2/A[7] ), 
        .D(n3685), .Y(n3980) );
  AOI22X1 U4233 ( .A(n4022), .B(\sub_x_1100_2/A[6] ), .C(n1819), .D(n2230), 
        .Y(n3983) );
  AOI22X1 U4234 ( .A(n1841), .B(n3496), .C(n3497), .D(n3910), .Y(n3993) );
  AOI22X1 U4235 ( .A(n4022), .B(\sub_x_1100_2/A[4] ), .C(n3721), .D(n2230), 
        .Y(n3982) );
  AOI22X1 U4236 ( .A(n2226), .B(\sub_x_1100_2/A[2] ), .C(n3722), .D(n2230), 
        .Y(n3959) );
  AOI22X1 U4237 ( .A(n1841), .B(n3654), .C(n2981), .D(n3910), .Y(n3960) );
  AOI22X1 U4238 ( .A(n2238), .B(n3498), .C(n2982), .D(n2251), .Y(n3961) );
  AOI22X1 U4239 ( .A(n2286), .B(n3495), .C(n2983), .D(n3908), .Y(n3962) );
  AOI22X1 U4240 ( .A(n2236), .B(n3361), .C(n2984), .D(n2239), .Y(n3964) );
  AOI22X1 U4241 ( .A(n2286), .B(n2907), .C(n3483), .D(n3908), .Y(n3992) );
  AOI22X1 U4242 ( .A(n2286), .B(n3968), .C(n4020), .D(n3908), .Y(n3998) );
  AOI22X1 U4243 ( .A(n2286), .B(n3292), .C(n3490), .D(n3908), .Y(n4004) );
  AOI22X1 U4244 ( .A(n2286), .B(n3294), .C(n3491), .D(n3908), .Y(n4008) );
  OR2X1 U4245 ( .A(n2286), .B(n3374), .Y(n4011) );
  OR2X1 U4246 ( .A(n2286), .B(n3375), .Y(n4014) );
  AOI22X1 U4247 ( .A(\ashr_1100_6/SH[1] ), .B(n3458), .C(n3461), .D(n3910), 
        .Y(n3999) );
  AOI22X1 U4248 ( .A(n1841), .B(n3493), .C(n3496), .D(n3910), .Y(n4005) );
  AOI22X1 U4249 ( .A(n1841), .B(n3497), .C(n3654), .D(n3910), .Y(n3984) );
  AOI22X1 U4250 ( .A(n2238), .B(n3500), .C(n2985), .D(n2251), .Y(n3985) );
  AOI22X1 U4251 ( .A(n2286), .B(n3482), .C(n2986), .D(n3908), .Y(n3987) );
  OAI21X1 U4252 ( .A(n3332), .B(n2239), .C(n2702), .Y(
        \arithmetic_logic_unit/N286 ) );
  AOI22X1 U4253 ( .A(n2238), .B(n3494), .C(n3498), .D(n2251), .Y(n3995) );
  AOI22X1 U4254 ( .A(n2286), .B(n3489), .C(n2987), .D(n3908), .Y(n3997) );
  OAI21X1 U4255 ( .A(n3333), .B(n2239), .C(n2703), .Y(
        \arithmetic_logic_unit/N288 ) );
  AOI22X1 U4256 ( .A(n2238), .B(n3467), .C(n3499), .D(n2251), .Y(n4001) );
  AOI22X1 U4257 ( .A(n2286), .B(n3280), .C(n2988), .D(n3908), .Y(n4003) );
  OAI21X1 U4258 ( .A(n3334), .B(n2239), .C(n2704), .Y(
        \arithmetic_logic_unit/N289 ) );
  NAND3X1 U4259 ( .A(memoryReadWrite), .B(n2221), .C(n4325), .Y(n4033) );
  NOR3X1 U4260 ( .A(n1001), .B(n4023), .C(n4029), .Y(n4363) );
  AOI22X1 U4261 ( .A(n1001), .B(memoryData[31]), .C(FRS2[31]), .D(n4023), .Y(
        n1354) );
  AOI22X1 U4262 ( .A(n1001), .B(memoryData[0]), .C(FRS2[0]), .D(n4023), .Y(
        n1352) );
  AOI22X1 U4263 ( .A(n1001), .B(memoryData[1]), .C(FRS2[1]), .D(n4023), .Y(
        n1350) );
  AOI22X1 U4264 ( .A(n1001), .B(memoryData[2]), .C(FRS2[2]), .D(n4023), .Y(
        n1348) );
  AOI22X1 U4265 ( .A(n1001), .B(memoryData[3]), .C(FRS2[3]), .D(n4023), .Y(
        n1346) );
  AOI22X1 U4266 ( .A(n1001), .B(memoryData[4]), .C(FRS2[4]), .D(n4023), .Y(
        n1344) );
  AOI22X1 U4267 ( .A(n1001), .B(memoryData[5]), .C(FRS2[5]), .D(n4023), .Y(
        n1342) );
  AOI22X1 U4268 ( .A(n1001), .B(memoryData[6]), .C(FRS2[6]), .D(n4023), .Y(
        n1340) );
  AOI22X1 U4269 ( .A(n1001), .B(memoryData[7]), .C(FRS2[7]), .D(n4023), .Y(
        n1338) );
  AOI22X1 U4270 ( .A(n1001), .B(memoryData[8]), .C(FRS2[8]), .D(n4023), .Y(
        n1336) );
  AOI22X1 U4271 ( .A(n1001), .B(memoryData[9]), .C(FRS2[9]), .D(n4023), .Y(
        n1334) );
  AOI22X1 U4272 ( .A(n1001), .B(memoryData[10]), .C(FRS2[10]), .D(n4023), .Y(
        n1332) );
  AOI22X1 U4273 ( .A(n1001), .B(memoryData[11]), .C(FRS2[11]), .D(n4023), .Y(
        n1330) );
  AOI22X1 U4274 ( .A(n1001), .B(memoryData[12]), .C(FRS2[12]), .D(n4023), .Y(
        n1328) );
  AOI22X1 U4275 ( .A(n1001), .B(memoryData[13]), .C(FRS2[13]), .D(n4023), .Y(
        n1326) );
  AOI22X1 U4276 ( .A(n1001), .B(memoryData[14]), .C(FRS2[14]), .D(n4023), .Y(
        n1324) );
  AOI22X1 U4277 ( .A(n1001), .B(memoryData[15]), .C(FRS2[15]), .D(n4023), .Y(
        n1322) );
  AOI22X1 U4278 ( .A(n1001), .B(memoryData[16]), .C(FRS2[16]), .D(n4023), .Y(
        n1320) );
  AOI22X1 U4279 ( .A(n1001), .B(memoryData[17]), .C(FRS2[17]), .D(n4023), .Y(
        n1318) );
  AOI22X1 U4280 ( .A(n1001), .B(memoryData[18]), .C(FRS2[18]), .D(n4023), .Y(
        n1316) );
  AOI22X1 U4281 ( .A(n1001), .B(memoryData[19]), .C(FRS2[19]), .D(n4023), .Y(
        n1314) );
  AOI22X1 U4282 ( .A(n1001), .B(memoryData[20]), .C(FRS2[20]), .D(n4023), .Y(
        n1312) );
  AOI22X1 U4283 ( .A(n1001), .B(memoryData[21]), .C(FRS2[21]), .D(n4023), .Y(
        n1310) );
  AOI22X1 U4284 ( .A(n1001), .B(memoryData[22]), .C(FRS2[22]), .D(n4023), .Y(
        n1308) );
  AOI22X1 U4285 ( .A(n1001), .B(memoryData[23]), .C(FRS2[23]), .D(n4023), .Y(
        n1306) );
  AOI22X1 U4286 ( .A(n1001), .B(memoryData[24]), .C(FRS2[24]), .D(n4023), .Y(
        n1304) );
  AOI22X1 U4287 ( .A(n1001), .B(memoryData[25]), .C(FRS2[25]), .D(n4023), .Y(
        n1302) );
  AOI22X1 U4288 ( .A(n1001), .B(memoryData[26]), .C(FRS2[26]), .D(n4023), .Y(
        n1300) );
  AOI22X1 U4289 ( .A(n1001), .B(memoryData[27]), .C(FRS2[27]), .D(n4023), .Y(
        n1298) );
  AOI22X1 U4290 ( .A(n1001), .B(memoryData[28]), .C(FRS2[28]), .D(n4023), .Y(
        n1296) );
  AOI22X1 U4291 ( .A(n1001), .B(memoryData[29]), .C(FRS2[29]), .D(n4023), .Y(
        n1294) );
  AOI22X1 U4292 ( .A(n1001), .B(memoryData[30]), .C(FRS2[30]), .D(n4023), .Y(
        n1289) );
  NAND3X1 U4293 ( .A(n2842), .B(n2927), .C(n2994), .Y(aluOperand1[31]) );
  NAND3X1 U4294 ( .A(n2844), .B(n2929), .C(n2996), .Y(aluOperand1[30]) );
  NAND3X1 U4295 ( .A(n2846), .B(n2931), .C(n2998), .Y(aluOperand1[29]) );
  NAND3X1 U4296 ( .A(n2848), .B(n2933), .C(n3000), .Y(aluOperand1[28]) );
  NAND3X1 U4297 ( .A(n2850), .B(n3632), .C(n3002), .Y(aluOperand1[27]) );
  AOI22X1 U4298 ( .A(n2266), .B(RS1[26]), .C(n2299), .D(pc[26]), .Y(n4037) );
  OAI21X1 U4299 ( .A(n4091), .B(n4038), .C(n2652), .Y(aluOperand1[26]) );
  AOI22X1 U4300 ( .A(n2266), .B(RS1[25]), .C(n2298), .D(pc[25]), .Y(n4039) );
  OAI21X1 U4301 ( .A(n4091), .B(n4040), .C(n2653), .Y(aluOperand1[25]) );
  AOI22X1 U4302 ( .A(n2266), .B(RS1[24]), .C(n2298), .D(pc[24]), .Y(n4041) );
  OAI21X1 U4303 ( .A(n4091), .B(n4042), .C(n2654), .Y(aluOperand1[24]) );
  AOI22X1 U4304 ( .A(n2266), .B(RS1[23]), .C(n2298), .D(pc[23]), .Y(n4043) );
  OAI21X1 U4305 ( .A(n4091), .B(n4044), .C(n2655), .Y(aluOperand1[23]) );
  AOI22X1 U4306 ( .A(n2266), .B(RS1[22]), .C(n2299), .D(pc[22]), .Y(n4045) );
  OAI21X1 U4307 ( .A(n4091), .B(n4046), .C(n2656), .Y(aluOperand1[22]) );
  AOI22X1 U4308 ( .A(n2266), .B(RS1[21]), .C(n2298), .D(pc[21]), .Y(n4047) );
  OAI21X1 U4309 ( .A(n4091), .B(n4048), .C(n2657), .Y(aluOperand1[21]) );
  AOI22X1 U4310 ( .A(n2266), .B(RS1[20]), .C(n2299), .D(pc[20]), .Y(n4049) );
  OAI21X1 U4311 ( .A(n4091), .B(n4050), .C(n2658), .Y(aluOperand1[20]) );
  AOI22X1 U4312 ( .A(n2266), .B(RS1[19]), .C(n2299), .D(pc[19]), .Y(n4051) );
  OAI21X1 U4313 ( .A(n4091), .B(n4052), .C(n2659), .Y(aluOperand1[19]) );
  AOI22X1 U4314 ( .A(n2266), .B(RS1[18]), .C(n2298), .D(pc[18]), .Y(n4053) );
  OAI21X1 U4315 ( .A(n4091), .B(n4054), .C(n2660), .Y(aluOperand1[18]) );
  AOI22X1 U4316 ( .A(n1833), .B(RS1[17]), .C(n2303), .D(pc[17]), .Y(n4055) );
  OAI21X1 U4317 ( .A(n4091), .B(n4056), .C(n2661), .Y(aluOperand1[17]) );
  AOI22X1 U4318 ( .A(n2266), .B(RS1[16]), .C(n2304), .D(pc[16]), .Y(n4057) );
  OAI21X1 U4319 ( .A(n4091), .B(n4058), .C(n2662), .Y(aluOperand1[16]) );
  AOI22X1 U4320 ( .A(RS1[15]), .B(n2278), .C(n2300), .D(pc[15]), .Y(n4059) );
  OAI21X1 U4321 ( .A(n4091), .B(n4060), .C(n2664), .Y(aluOperand1[15]) );
  AOI22X1 U4322 ( .A(n3696), .B(RS1[14]), .C(n2301), .D(pc[14]), .Y(n4061) );
  OAI21X1 U4323 ( .A(n4091), .B(n4062), .C(n2380), .Y(aluOperand1[14]) );
  AOI22X1 U4324 ( .A(n1832), .B(RS1[13]), .C(n2304), .D(pc[13]), .Y(n4063) );
  OAI21X1 U4325 ( .A(n4091), .B(n4064), .C(n2666), .Y(aluOperand1[13]) );
  AOI22X1 U4326 ( .A(n1813), .B(RS1[12]), .C(n2304), .D(pc[12]), .Y(n4065) );
  OAI21X1 U4327 ( .A(n4091), .B(n4066), .C(n2668), .Y(aluOperand1[12]) );
  AOI22X1 U4328 ( .A(n1813), .B(RS1[11]), .C(n2302), .D(pc[11]), .Y(n4067) );
  OAI21X1 U4329 ( .A(n4091), .B(n4068), .C(n2669), .Y(aluOperand1[11]) );
  AOI22X1 U4330 ( .A(RS1[10]), .B(n3697), .C(n2237), .D(pc[10]), .Y(n4069) );
  OAI21X1 U4331 ( .A(n4091), .B(n4070), .C(n2381), .Y(aluOperand1[10]) );
  AOI22X1 U4332 ( .A(n3700), .B(RS1[9]), .C(n2301), .D(pc[9]), .Y(n4071) );
  AOI22X1 U4333 ( .A(n4089), .B(RS1[8]), .C(n2303), .D(pc[8]), .Y(n4073) );
  OAI21X1 U4334 ( .A(n4091), .B(n4074), .C(n2670), .Y(aluOperand1[8]) );
  AOI22X1 U4335 ( .A(n4089), .B(RS1[7]), .C(n2300), .D(pc[7]), .Y(n4075) );
  OAI21X1 U4336 ( .A(n4091), .B(n4076), .C(n2672), .Y(aluOperand1[7]) );
  AOI22X1 U4337 ( .A(n3699), .B(RS1[6]), .C(n2302), .D(pc[6]), .Y(n4077) );
  OAI21X1 U4338 ( .A(n4091), .B(n4078), .C(n2674), .Y(aluOperand1[6]) );
  AOI22X1 U4339 ( .A(n4089), .B(RS1[5]), .C(n2237), .D(pc[5]), .Y(n4079) );
  OAI21X1 U4340 ( .A(n4091), .B(n4080), .C(n2675), .Y(aluOperand1[5]) );
  AOI22X1 U4341 ( .A(n3695), .B(RS1[4]), .C(n2300), .D(pc[4]), .Y(n4081) );
  OAI21X1 U4342 ( .A(n4091), .B(n4082), .C(n2677), .Y(aluOperand1[4]) );
  AOI22X1 U4343 ( .A(n3698), .B(RS1[3]), .C(n2301), .D(pc[3]), .Y(n4083) );
  OAI21X1 U4344 ( .A(n4091), .B(n4084), .C(n2678), .Y(aluOperand1[3]) );
  AOI22X1 U4345 ( .A(RS1[2]), .B(n3701), .C(n2302), .D(pc[2]), .Y(n4085) );
  OAI21X1 U4346 ( .A(n4091), .B(n4086), .C(n2679), .Y(aluOperand1[2]) );
  AOI22X1 U4347 ( .A(RS1[1]), .B(n4089), .C(n2302), .D(pc[1]), .Y(n4087) );
  OAI21X1 U4348 ( .A(n4091), .B(n4088), .C(n2680), .Y(aluOperand1[1]) );
  OAI21X1 U4349 ( .A(n4091), .B(n4090), .C(n2383), .Y(aluOperand1[0]) );
  AOI22X1 U4350 ( .A(n2282), .B(RS2[31]), .C(n2306), .D(immediate[31]), .Y(
        n4292) );
  AOI22X1 U4351 ( .A(n2282), .B(RS2[30]), .C(n2306), .D(immediate[30]), .Y(
        n4291) );
  AOI22X1 U4352 ( .A(n2282), .B(RS2[29]), .C(n2306), .D(immediate[29]), .Y(
        n4290) );
  AOI22X1 U4353 ( .A(n2282), .B(RS2[28]), .C(n2306), .D(immediate[28]), .Y(
        n4286) );
  AOI22X1 U4354 ( .A(n2281), .B(RS2[27]), .C(n2306), .D(immediate[27]), .Y(
        n4279) );
  AOI22X1 U4355 ( .A(n2282), .B(RS2[26]), .C(n2306), .D(immediate[26]), .Y(
        n4268) );
  AOI22X1 U4356 ( .A(n2281), .B(RS2[25]), .C(n2306), .D(immediate[25]), .Y(
        n4261) );
  AOI22X1 U4357 ( .A(n2282), .B(RS2[24]), .C(n2306), .D(immediate[24]), .Y(
        n4253) );
  AOI22X1 U4358 ( .A(n2282), .B(RS2[23]), .C(n2306), .D(immediate[23]), .Y(
        n4246) );
  AOI22X1 U4359 ( .A(n2282), .B(RS2[22]), .C(n2306), .D(immediate[22]), .Y(
        n4238) );
  AOI22X1 U4360 ( .A(n2282), .B(RS2[21]), .C(n2306), .D(immediate[21]), .Y(
        n4230) );
  AOI22X1 U4361 ( .A(n2281), .B(RS2[20]), .C(n2306), .D(immediate[20]), .Y(
        n4229) );
  AOI22X1 U4362 ( .A(n2282), .B(RS2[19]), .C(n2306), .D(immediate[19]), .Y(
        n4228) );
  AOI22X1 U4363 ( .A(n2265), .B(RS2[17]), .C(n2306), .D(immediate[17]), .Y(
        n4221) );
  AOI22X1 U4364 ( .A(n2242), .B(RS2[16]), .C(n2306), .D(immediate[16]), .Y(
        n4093) );
  AOI22X1 U4365 ( .A(n2215), .B(RS2[15]), .C(n4102), .D(immediate[15]), .Y(
        n4215) );
  AOI22X1 U4366 ( .A(n2215), .B(RS2[14]), .C(n4102), .D(immediate[14]), .Y(
        n4214) );
  AOI22X1 U4367 ( .A(n2216), .B(RS2[13]), .C(n4102), .D(immediate[13]), .Y(
        n4213) );
  AOI22X1 U4368 ( .A(n2216), .B(RS2[12]), .C(n4102), .D(immediate[12]), .Y(
        n4212) );
  AOI22X1 U4369 ( .A(n2216), .B(RS2[11]), .C(n4102), .D(immediate[11]), .Y(
        n4205) );
  AOI22X1 U4370 ( .A(n2215), .B(RS2[10]), .C(n4102), .D(immediate[10]), .Y(
        n4094) );
  AOI22X1 U4371 ( .A(n2280), .B(RS2[9]), .C(n4102), .D(immediate[9]), .Y(n4095) );
  AOI22X1 U4372 ( .A(n2216), .B(RS2[8]), .C(n4102), .D(immediate[8]), .Y(n4096) );
  AOI22X1 U4373 ( .A(n2215), .B(RS2[7]), .C(n4102), .D(immediate[7]), .Y(n4097) );
  AOI22X1 U4374 ( .A(n2280), .B(RS2[6]), .C(n4102), .D(immediate[6]), .Y(n4098) );
  AOI22X1 U4375 ( .A(n2280), .B(RS2[5]), .C(n4102), .D(immediate[5]), .Y(n4099) );
  AOI22X1 U4376 ( .A(n2216), .B(RS2[4]), .C(n4102), .D(immediate[4]), .Y(n4194) );
  AOI22X1 U4377 ( .A(n1830), .B(n4100), .C(n2280), .D(RS2[2]), .Y(n4101) );
  NOR3X1 U4378 ( .A(n4369), .B(n4368), .C(n2432), .Y(n4293) );
  NOR3X1 U4379 ( .A(n2272), .B(n4329), .C(n2404), .Y(n4332) );
  AOI21X1 U4380 ( .A(n4115), .B(n2355), .C(n4332), .Y(n4106) );
  NAND3X1 U4381 ( .A(n3720), .B(n2290), .C(n4107), .Y(n4165) );
  NAND3X1 U4382 ( .A(n3719), .B(n2267), .C(n4108), .Y(n4146) );
  OAI21X1 U4383 ( .A(n3378), .B(n2402), .C(n4325), .Y(n4109) );
  AOI21X1 U4384 ( .A(n4332), .B(n4325), .C(n4136), .Y(n4140) );
  AOI21X1 U4385 ( .A(n2220), .B(\funct3[0] ), .C(funct3[1]), .Y(n4150) );
  MUX2X1 U4386 ( .B(n2883), .A(n4110), .S(n4334), .Y(n4111) );
  NOR3X1 U4387 ( .A(n3555), .B(n4112), .C(n4111), .Y(n4362) );
  NAND3X1 U4388 ( .A(n4120), .B(n4113), .C(n3506), .Y(n4114) );
  NAND3X1 U4389 ( .A(n3673), .B(n2922), .C(n3004), .Y(n4116) );
  MUX2X1 U4390 ( .B(n2887), .A(n1145), .S(aluZeroRegister), .Y(n4118) );
  OAI21X1 U4391 ( .A(n3653), .B(n4118), .C(n4334), .Y(n4119) );
  MUX2X1 U4392 ( .B(n2885), .A(n2914), .S(n4120), .Y(n4121) );
  AOI22X1 U4393 ( .A(n2920), .B(n4121), .C(n3318), .D(n2990), .Y(n504) );
  AOI22X1 U4394 ( .A(n3674), .B(n4122), .C(n3724), .D(n2362), .Y(n4127) );
  MUX2X1 U4395 ( .B(n1145), .A(n2454), .S(aluZeroRegister), .Y(n4123) );
  AOI21X1 U4396 ( .A(aluSignRegister), .B(n2220), .C(n4123), .Y(n4124) );
  OAI21X1 U4397 ( .A(n2879), .B(n2309), .C(n4336), .Y(n4125) );
  AOI21X1 U4398 ( .A(n3719), .B(n4330), .C(n2437), .Y(n4133) );
  AOI21X1 U4399 ( .A(n4334), .B(n4125), .C(n3304), .Y(n4126) );
  AOI21X1 U4400 ( .A(memoryReady), .B(n4336), .C(n61), .Y(n4132) );
  AOI21X1 U4401 ( .A(memoryReady), .B(n4334), .C(n3724), .Y(n4128) );
  MUX2X1 U4402 ( .B(n3674), .A(n2913), .S(n4366), .Y(n4129) );
  NAND3X1 U4403 ( .A(n3187), .B(n4131), .C(n2309), .Y(n4144) );
  AOI21X1 U4404 ( .A(n4168), .B(n2353), .C(n3554), .Y(n4134) );
  NOR3X1 U4405 ( .A(n3039), .B(n3042), .C(n3046), .Y(n515) );
  OAI21X1 U4406 ( .A(n4168), .B(n3506), .C(n3726), .Y(n517) );
  NOR3X1 U4407 ( .A(n3726), .B(n4365), .C(n2269), .Y(n4337) );
  NOR3X1 U4408 ( .A(n2219), .B(n3555), .C(n2471), .Y(n518) );
  NOR3X1 U4409 ( .A(n2467), .B(n4333), .C(n2362), .Y(n4142) );
  NOR3X1 U4410 ( .A(n3548), .B(n3553), .C(n2475), .Y(n4135) );
  NOR3X1 U4411 ( .A(n3040), .B(n2475), .C(n3554), .Y(n526) );
  NAND3X1 U4412 ( .A(n2270), .B(n2354), .C(n3007), .Y(n4138) );
  NAND3X1 U4413 ( .A(n4136), .B(n2309), .C(n3673), .Y(n4137) );
  AOI21X1 U4414 ( .A(n4168), .B(n2854), .C(n2800), .Y(n533) );
  NAND3X1 U4415 ( .A(n3549), .B(n2365), .C(n4139), .Y(n4141) );
  AOI22X1 U4416 ( .A(n3548), .B(n2919), .C(n3726), .D(n3552), .Y(n4143) );
  NOR3X1 U4417 ( .A(n2360), .B(n2367), .C(n2288), .Y(n4361) );
  OAI21X1 U4418 ( .A(n4365), .B(n4366), .C(n4334), .Y(n535) );
  OAI21X1 U4419 ( .A(n4334), .B(n4366), .C(n4365), .Y(n543) );
  NOR3X1 U4420 ( .A(n4337), .B(n3554), .C(n3048), .Y(n544) );
  NOR3X1 U4421 ( .A(n3726), .B(n2212), .C(n3725), .Y(n4166) );
  NOR3X1 U4422 ( .A(n4166), .B(n3674), .C(n2449), .Y(n547) );
  AOI22X1 U4423 ( .A(n4168), .B(n3378), .C(n3186), .D(n4145), .Y(n549) );
  NOR3X1 U4424 ( .A(n2279), .B(n2221), .C(n3562), .Y(n4161) );
  NAND3X1 U4425 ( .A(n4151), .B(n4168), .C(n3008), .Y(n551) );
  NOR3X1 U4426 ( .A(n3503), .B(n4159), .C(n3052), .Y(n4149) );
  OAI21X1 U4427 ( .A(n4149), .B(n3376), .C(n4161), .Y(n4154) );
  NAND3X1 U4428 ( .A(n3376), .B(n4163), .C(n4151), .Y(n4152) );
  NAND3X1 U4429 ( .A(n4154), .B(n4153), .C(n2992), .Y(n4156) );
  AOI21X1 U4430 ( .A(n4168), .B(n2855), .C(n4155), .Y(n4360) );
  NAND3X1 U4431 ( .A(n4168), .B(n138), .C(n3321), .Y(n4157) );
  AOI21X1 U4432 ( .A(n1144), .B(n3253), .C(n2801), .Y(n4158) );
  NAND3X1 U4433 ( .A(n3254), .B(n4168), .C(n3010), .Y(n555) );
  AOI21X1 U4434 ( .A(n3517), .B(n4160), .C(n1138), .Y(n4162) );
  OAI21X1 U4435 ( .A(n3503), .B(n2960), .C(n4161), .Y(n4164) );
  NAND3X1 U4436 ( .A(n3719), .B(n4164), .C(n3012), .Y(n4167) );
  AOI21X1 U4437 ( .A(n4168), .B(n2856), .C(n4166), .Y(n557) );
  AOI22X1 U4438 ( .A(n4371), .B(ir[20]), .C(ir_7), .D(n4370), .Y(n4169) );
  MUX2X1 U4439 ( .B(ir[21]), .A(ir_8), .S(instructionType[1]), .Y(n4170) );
  MUX2X1 U4440 ( .B(ir[22]), .A(ir_9), .S(instructionType[1]), .Y(n4171) );
  MUX2X1 U4441 ( .B(ir[23]), .A(ir_10), .S(instructionType[1]), .Y(n4172) );
  MUX2X1 U4442 ( .B(ir[24]), .A(ir_11), .S(instructionType[1]), .Y(n4174) );
  NAND3X1 U4443 ( .A(instructionType[2]), .B(n2935), .C(n4175), .Y(n4180) );
  NAND3X1 U4444 ( .A(instructionType[0]), .B(n4372), .C(n3014), .Y(n4179) );
  OAI21X1 U4445 ( .A(instructionType[0]), .B(funct7[6]), .C(n3723), .Y(n4176)
         );
  AOI21X1 U4446 ( .A(n4371), .B(n4177), .C(n4176), .Y(n4178) );
  OAI21X1 U4447 ( .A(\funct3[0] ), .B(n4372), .C(n4181), .Y(n871) );
  OAI21X1 U4448 ( .A(funct3[1]), .B(n4372), .C(n4181), .Y(n873) );
  OAI21X1 U4449 ( .A(n2220), .B(n4372), .C(n4181), .Y(n875) );
  OAI21X1 U4450 ( .A(ir[15]), .B(n4372), .C(n4181), .Y(n877) );
  OAI21X1 U4451 ( .A(ir[16]), .B(n4372), .C(n4181), .Y(n879) );
  OAI21X1 U4452 ( .A(n4372), .B(ir[17]), .C(n4181), .Y(n881) );
  OAI21X1 U4453 ( .A(n4372), .B(ir[18]), .C(n4181), .Y(n883) );
  OAI21X1 U4454 ( .A(n4372), .B(ir[19]), .C(n4181), .Y(n885) );
  OAI21X1 U4455 ( .A(ir[20]), .B(n3723), .C(n3677), .Y(n887) );
  OAI21X1 U4456 ( .A(ir[21]), .B(n3723), .C(n3677), .Y(n889) );
  OAI21X1 U4457 ( .A(ir[22]), .B(n3723), .C(n3677), .Y(n891) );
  OAI21X1 U4458 ( .A(ir[23]), .B(n3723), .C(n3677), .Y(n893) );
  OAI21X1 U4459 ( .A(ir[24]), .B(n3723), .C(n3677), .Y(n895) );
  OAI21X1 U4460 ( .A(funct7[0]), .B(n3723), .C(n3677), .Y(n897) );
  OAI21X1 U4461 ( .A(funct7[1]), .B(n3723), .C(n3677), .Y(n899) );
  OAI21X1 U4462 ( .A(funct7[2]), .B(n3723), .C(n3677), .Y(n901) );
  OAI21X1 U4463 ( .A(funct7[3]), .B(n3723), .C(n3677), .Y(n903) );
  OAI21X1 U4464 ( .A(funct7[4]), .B(n3723), .C(n3677), .Y(n905) );
  OAI21X1 U4465 ( .A(funct7[5]), .B(n3723), .C(n3677), .Y(n907) );
  AOI21X1 U4466 ( .A(n3704), .B(n3910), .C(n3709), .Y(n4184) );
  MUX2X1 U4467 ( .B(n2241), .A(n4269), .S(n3722), .Y(n4182) );
  OAI21X1 U4468 ( .A(n4182), .B(n3709), .C(n1841), .Y(n4183) );
  OAI21X1 U4469 ( .A(n3758), .B(n2961), .C(n4183), .Y(n4185) );
  AOI21X1 U4470 ( .A(\arithmetic_logic_unit/N90 ), .B(n4026), .C(n4185), .Y(
        n4186) );
  NAND3X1 U4471 ( .A(n2830), .B(n2398), .C(n3016), .Y(n4187) );
  AOI21X1 U4472 ( .A(\arithmetic_logic_unit/N284 ), .B(aluOperation[3]), .C(
        n2802), .Y(n913) );
  AOI21X1 U4473 ( .A(n3704), .B(n3712), .C(n3709), .Y(n4190) );
  MUX2X1 U4474 ( .B(n2241), .A(n4269), .S(n3721), .Y(n4188) );
  OAI21X1 U4475 ( .A(n4188), .B(n3709), .C(n2286), .Y(n4189) );
  OAI21X1 U4476 ( .A(n3750), .B(n2962), .C(n4189), .Y(n4191) );
  AOI21X1 U4477 ( .A(\arithmetic_logic_unit/N92 ), .B(n4026), .C(n4191), .Y(
        n4192) );
  NAND3X1 U4478 ( .A(n2831), .B(n2400), .C(n2369), .Y(n4193) );
  AOI21X1 U4479 ( .A(\arithmetic_logic_unit/N286 ), .B(aluOperation[3]), .C(
        n2803), .Y(n917) );
  MUX2X1 U4480 ( .B(n3704), .A(n1381), .S(n1819), .Y(n4195) );
  OAI21X1 U4481 ( .A(n2241), .B(n1831), .C(n2240), .Y(n4196) );
  AOI22X1 U4482 ( .A(n1831), .B(n2909), .C(n1819), .D(n4196), .Y(n4197) );
  AOI21X1 U4483 ( .A(\arithmetic_logic_unit/N288 ), .B(aluOperation[3]), .C(
        n2822), .Y(n4199) );
  AOI22X1 U4484 ( .A(n4293), .B(n2901), .C(n4027), .D(
        \arithmetic_logic_unit/N126 ), .Y(n4198) );
  MUX2X1 U4485 ( .B(n3704), .A(n1381), .S(\sub_x_1100_2/A[6] ), .Y(n4200) );
  OAI21X1 U4486 ( .A(n2241), .B(n2292), .C(n2240), .Y(n4201) );
  AOI22X1 U4487 ( .A(n2292), .B(n2911), .C(\sub_x_1100_2/A[6] ), .D(n4201), 
        .Y(n4202) );
  AOI21X1 U4488 ( .A(\arithmetic_logic_unit/N289 ), .B(aluOperation[3]), .C(
        n2824), .Y(n4204) );
  AOI22X1 U4489 ( .A(n4293), .B(n2903), .C(n4027), .D(
        \arithmetic_logic_unit/N127 ), .Y(n4203) );
  AOI21X1 U4490 ( .A(n3704), .B(n3252), .C(n3709), .Y(n4208) );
  MUX2X1 U4491 ( .B(n2241), .A(n4269), .S(\sub_x_1100_2/A[11] ), .Y(n4206) );
  OAI21X1 U4492 ( .A(n4206), .B(n3709), .C(\lt_x_1100_4/B[11] ), .Y(n4207) );
  OAI21X1 U4493 ( .A(n3764), .B(n2963), .C(n4207), .Y(n4209) );
  AOI21X1 U4494 ( .A(n4293), .B(n2392), .C(n4209), .Y(n4210) );
  NAND3X1 U4495 ( .A(n2389), .B(n2937), .C(n3018), .Y(n4211) );
  AOI21X1 U4496 ( .A(\arithmetic_logic_unit/N132 ), .B(n4027), .C(n2804), .Y(
        n933) );
  AOI21X1 U4497 ( .A(n3704), .B(n1827), .C(n3709), .Y(n4218) );
  MUX2X1 U4498 ( .B(n2241), .A(n4269), .S(n2060), .Y(n4216) );
  OAI21X1 U4499 ( .A(n4216), .B(n3709), .C(\lt_x_1100_4/B[15] ), .Y(n4217) );
  OAI21X1 U4500 ( .A(n3762), .B(n2964), .C(n4217), .Y(n4219) );
  AOI21X1 U4501 ( .A(\arithmetic_logic_unit/N266 ), .B(n4293), .C(n4219), .Y(
        n4220) );
  AOI21X1 U4502 ( .A(\arithmetic_logic_unit/N136 ), .B(n4027), .C(n2310), .Y(
        n941) );
  AOI21X1 U4503 ( .A(n3704), .B(n3248), .C(n3709), .Y(n4224) );
  MUX2X1 U4504 ( .B(n2241), .A(n4269), .S(aluOperand1[17]), .Y(n4222) );
  OAI21X1 U4505 ( .A(n4222), .B(n3709), .C(\lt_x_1100_4/B[17] ), .Y(n4223) );
  OAI21X1 U4506 ( .A(n3761), .B(n2965), .C(n4223), .Y(n4225) );
  AOI21X1 U4507 ( .A(\arithmetic_logic_unit/N300 ), .B(aluOperation[3]), .C(
        n4225), .Y(n4226) );
  NAND3X1 U4508 ( .A(n2832), .B(n2940), .C(n3021), .Y(n4227) );
  AOI21X1 U4509 ( .A(\arithmetic_logic_unit/N138 ), .B(n4027), .C(n2806), .Y(
        n945) );
  AOI21X1 U4510 ( .A(n3704), .B(n3245), .C(n3709), .Y(n4233) );
  MUX2X1 U4511 ( .B(n2241), .A(n4269), .S(aluOperand1[21]), .Y(n4231) );
  OAI21X1 U4512 ( .A(n4231), .B(n3709), .C(\lt_x_1100_4/B[21] ), .Y(n4232) );
  OAI21X1 U4513 ( .A(n4234), .B(n2966), .C(n4232), .Y(n4235) );
  AOI21X1 U4514 ( .A(aluOperation[3]), .B(n2441), .C(n4235), .Y(n4236) );
  NAND3X1 U4515 ( .A(n2833), .B(n2942), .C(n3023), .Y(n4237) );
  AOI21X1 U4516 ( .A(\arithmetic_logic_unit/N142 ), .B(n4027), .C(n2807), .Y(
        n953) );
  AOI21X1 U4517 ( .A(n3704), .B(n3244), .C(n3709), .Y(n4241) );
  MUX2X1 U4518 ( .B(n2241), .A(n4269), .S(aluOperand1[22]), .Y(n4239) );
  OAI21X1 U4519 ( .A(n4239), .B(n3709), .C(\lt_x_1100_4/B[22] ), .Y(n4240) );
  OAI21X1 U4520 ( .A(n4242), .B(n2967), .C(n4240), .Y(n4243) );
  AOI21X1 U4521 ( .A(aluOperation[3]), .B(n2443), .C(n4243), .Y(n4244) );
  NAND3X1 U4522 ( .A(n2834), .B(n2944), .C(n3025), .Y(n4245) );
  AOI21X1 U4523 ( .A(\arithmetic_logic_unit/N143 ), .B(n4027), .C(n2808), .Y(
        n955) );
  AOI21X1 U4524 ( .A(n3704), .B(n3243), .C(n3709), .Y(n4249) );
  MUX2X1 U4525 ( .B(n2241), .A(n4269), .S(aluOperand1[23]), .Y(n4247) );
  OAI21X1 U4526 ( .A(n4247), .B(n3709), .C(\lt_x_1100_4/B[23] ), .Y(n4248) );
  OAI21X1 U4527 ( .A(n3757), .B(n2968), .C(n4248), .Y(n4250) );
  AOI21X1 U4528 ( .A(aluOperation[3]), .B(n2445), .C(n4250), .Y(n4251) );
  NAND3X1 U4529 ( .A(n2835), .B(n2946), .C(n3027), .Y(n4252) );
  AOI21X1 U4530 ( .A(\arithmetic_logic_unit/N144 ), .B(n4027), .C(n2809), .Y(
        n957) );
  AOI21X1 U4531 ( .A(n3704), .B(n3242), .C(n3709), .Y(n4256) );
  MUX2X1 U4532 ( .B(n2241), .A(n4269), .S(aluOperand1[24]), .Y(n4254) );
  OAI21X1 U4533 ( .A(n4254), .B(n3709), .C(\lt_x_1100_4/B[24] ), .Y(n4255) );
  OAI21X1 U4534 ( .A(n4257), .B(n2969), .C(n4255), .Y(n4258) );
  AOI21X1 U4535 ( .A(aluOperation[3]), .B(n2860), .C(n4258), .Y(n4259) );
  NAND3X1 U4536 ( .A(n2836), .B(n2948), .C(n3029), .Y(n4260) );
  AOI21X1 U4537 ( .A(\arithmetic_logic_unit/N145 ), .B(n4027), .C(n2810), .Y(
        n959) );
  AOI21X1 U4538 ( .A(n3704), .B(n3241), .C(n3709), .Y(n4264) );
  MUX2X1 U4539 ( .B(n2241), .A(n4269), .S(aluOperand1[25]), .Y(n4262) );
  OAI21X1 U4540 ( .A(n4262), .B(n3709), .C(\lt_x_1100_4/B[25] ), .Y(n4263) );
  OAI21X1 U4541 ( .A(n3756), .B(n2970), .C(n4263), .Y(n4265) );
  AOI21X1 U4542 ( .A(aluOperation[3]), .B(n2862), .C(n4265), .Y(n4266) );
  NAND3X1 U4543 ( .A(n2837), .B(n2950), .C(n3031), .Y(n4267) );
  AOI21X1 U4544 ( .A(\arithmetic_logic_unit/N146 ), .B(n4027), .C(n2811), .Y(
        n961) );
  AOI21X1 U4545 ( .A(n3704), .B(n3240), .C(n3709), .Y(n4272) );
  MUX2X1 U4546 ( .B(n2241), .A(n4269), .S(aluOperand1[26]), .Y(n4270) );
  OAI21X1 U4547 ( .A(n4270), .B(n3709), .C(\lt_x_1100_4/B[26] ), .Y(n4271) );
  OAI21X1 U4548 ( .A(n3755), .B(n2971), .C(n4271), .Y(n4273) );
  AOI21X1 U4549 ( .A(aluOperation[3]), .B(n2864), .C(n4273), .Y(n4274) );
  NAND3X1 U4550 ( .A(n2838), .B(n2952), .C(n3033), .Y(n4275) );
  AOI21X1 U4551 ( .A(\arithmetic_logic_unit/N147 ), .B(n4027), .C(n2812), .Y(
        n963) );
  OAI21X1 U4552 ( .A(n2241), .B(\sub_x_1100_2/A[27] ), .C(n2240), .Y(n4276) );
  AOI21X1 U4553 ( .A(n1381), .B(\sub_x_1100_2/A[27] ), .C(n4276), .Y(n4278) );
  OAI21X1 U4554 ( .A(n2241), .B(\lt_x_1100_4/B[27] ), .C(n2240), .Y(n4277) );
  OAI21X1 U4555 ( .A(n3258), .B(n2972), .C(n2705), .Y(n4280) );
  AOI21X1 U4556 ( .A(aluOperation[3]), .B(n2866), .C(n4280), .Y(n4281) );
  NAND3X1 U4557 ( .A(n2839), .B(n2954), .C(n3035), .Y(n4282) );
  AOI21X1 U4558 ( .A(\arithmetic_logic_unit/N148 ), .B(n4027), .C(n2813), .Y(
        n965) );
  OAI21X1 U4559 ( .A(n2241), .B(\sub_x_1100_2/A[28] ), .C(n2240), .Y(n4283) );
  AOI21X1 U4560 ( .A(n1381), .B(\sub_x_1100_2/A[28] ), .C(n4283), .Y(n4285) );
  OAI21X1 U4561 ( .A(n2241), .B(\lt_x_1100_4/B[28] ), .C(n2240), .Y(n4284) );
  OAI21X1 U4562 ( .A(n3257), .B(n2973), .C(n2707), .Y(n4287) );
  AOI21X1 U4563 ( .A(aluOperation[3]), .B(n2868), .C(n4287), .Y(n4288) );
  NAND3X1 U4564 ( .A(n2840), .B(n2956), .C(n2371), .Y(n4289) );
  AOI21X1 U4565 ( .A(\arithmetic_logic_unit/N117 ), .B(n4026), .C(n2815), .Y(
        n967) );
  AOI22X1 U4566 ( .A(n4028), .B(pc[2]), .C(n4340), .D(aluResult[2]), .Y(n4294)
         );
  AOI22X1 U4567 ( .A(n4028), .B(pc[10]), .C(n4340), .D(aluResult[10]), .Y(
        n4295) );
  AOI22X1 U4568 ( .A(n4028), .B(pc[11]), .C(n4340), .D(aluResult[11]), .Y(
        n4296) );
  AOI22X1 U4569 ( .A(n4028), .B(pc[12]), .C(n4340), .D(aluResult[12]), .Y(
        n4297) );
  AOI22X1 U4570 ( .A(n4028), .B(pc[13]), .C(n4340), .D(aluResult[13]), .Y(
        n4298) );
  AOI22X1 U4571 ( .A(n4028), .B(pc[14]), .C(n4340), .D(aluResult[14]), .Y(
        n4299) );
  AOI22X1 U4572 ( .A(n4028), .B(pc[15]), .C(n4340), .D(aluResult[15]), .Y(
        n4300) );
  AOI22X1 U4573 ( .A(n4028), .B(pc[17]), .C(n4340), .D(aluResult[17]), .Y(
        n4301) );
  AOI22X1 U4574 ( .A(n4028), .B(pc[18]), .C(n4340), .D(aluResult[18]), .Y(
        n4302) );
  AOI22X1 U4575 ( .A(n4028), .B(pc[19]), .C(n4340), .D(aluResult[19]), .Y(
        n4303) );
  AOI22X1 U4576 ( .A(n4028), .B(pc[1]), .C(n4340), .D(aluResult[1]), .Y(n4304)
         );
  AOI22X1 U4577 ( .A(n4028), .B(pc[20]), .C(n4340), .D(aluResult[20]), .Y(
        n4305) );
  AOI22X1 U4578 ( .A(n4028), .B(pc[21]), .C(n4340), .D(aluResult[21]), .Y(
        n4306) );
  AOI22X1 U4579 ( .A(n4028), .B(pc[22]), .C(n4340), .D(aluResult[22]), .Y(
        n4307) );
  AOI22X1 U4580 ( .A(n4028), .B(pc[23]), .C(n4340), .D(aluResult[23]), .Y(
        n4308) );
  AOI22X1 U4581 ( .A(n4028), .B(pc[24]), .C(n4340), .D(aluResult[24]), .Y(
        n4309) );
  AOI22X1 U4582 ( .A(n4028), .B(pc[25]), .C(n4340), .D(aluResult[25]), .Y(
        n4310) );
  AOI22X1 U4583 ( .A(n4028), .B(pc[26]), .C(n4340), .D(aluResult[26]), .Y(
        n4311) );
  AOI22X1 U4584 ( .A(n4028), .B(pc[27]), .C(n4340), .D(aluResult[27]), .Y(
        n4312) );
  AOI22X1 U4585 ( .A(n4028), .B(pc[29]), .C(n4340), .D(aluResult[29]), .Y(
        n4313) );
  AOI22X1 U4586 ( .A(n4028), .B(pc[3]), .C(n4340), .D(aluResult[3]), .Y(n4314)
         );
  AOI22X1 U4587 ( .A(n4028), .B(pc[4]), .C(n4340), .D(aluResult[4]), .Y(n4315)
         );
  AOI22X1 U4588 ( .A(n4028), .B(pc[5]), .C(n4340), .D(aluResult[5]), .Y(n4316)
         );
  AOI22X1 U4589 ( .A(n4028), .B(pc[6]), .C(n4340), .D(aluResult[6]), .Y(n4317)
         );
  AOI22X1 U4590 ( .A(n4028), .B(pc[7]), .C(n4340), .D(aluResult[7]), .Y(n4318)
         );
  AOI22X1 U4591 ( .A(n4028), .B(pc[9]), .C(n4340), .D(aluResult[9]), .Y(n4319)
         );
  NAND3X1 U4592 ( .A(n4325), .B(n2923), .C(n4320), .Y(n4321) );
  NOR3X1 U4593 ( .A(n2358), .B(n3558), .C(n3045), .Y(n4359) );
  MUX2X1 U4594 ( .B(n1851), .A(n3720), .S(n2279), .Y(n4323) );
  OAI21X1 U4595 ( .A(opcode[5]), .B(n2222), .C(n3546), .Y(n4324) );
  AOI21X1 U4596 ( .A(n4326), .B(n2405), .C(n3718), .Y(N466) );
  NAND3X1 U4597 ( .A(opcode[5]), .B(n3720), .C(n2290), .Y(n4327) );
  AOI21X1 U4598 ( .A(n1851), .B(n4329), .C(n2826), .Y(n4331) );
  OAI21X1 U4599 ( .A(n3546), .B(n2405), .C(n2709), .Y(N467) );
  AOI21X1 U4600 ( .A(n3725), .B(n3674), .C(n2362), .Y(n4335) );
  OAI21X1 U4601 ( .A(n3724), .B(n2309), .C(n4336), .Y(n4338) );
  AOI21X1 U4602 ( .A(n3726), .B(n4338), .C(n4337), .Y(n4339) );
  AOI21X1 U4603 ( .A(n3155), .B(n2857), .C(n3558), .Y(N924) );
  AOI22X1 U4604 ( .A(n4028), .B(pc[0]), .C(n4340), .D(aluResult[0]), .Y(n4341)
         );
  AOI22X1 U4605 ( .A(n4090), .B(instructionOrData), .C(n1034), .D(n4342), .Y(
        memoryAddress[0]) );
  AOI22X1 U4606 ( .A(n4088), .B(instructionOrData), .C(n1034), .D(n4343), .Y(
        memoryAddress[1]) );
  AOI22X1 U4607 ( .A(n4086), .B(instructionOrData), .C(n1034), .D(n4344), .Y(
        memoryAddress[2]) );
  AOI22X1 U4608 ( .A(n4084), .B(instructionOrData), .C(n1034), .D(n4345), .Y(
        memoryAddress[3]) );
  AOI22X1 U4609 ( .A(n4082), .B(instructionOrData), .C(n1034), .D(n4346), .Y(
        memoryAddress[4]) );
  AOI22X1 U4610 ( .A(n4080), .B(instructionOrData), .C(n1034), .D(n4347), .Y(
        memoryAddress[5]) );
  AOI22X1 U4611 ( .A(n4078), .B(instructionOrData), .C(n1034), .D(n4348), .Y(
        memoryAddress[6]) );
  AOI22X1 U4612 ( .A(n4076), .B(instructionOrData), .C(n1034), .D(n4349), .Y(
        memoryAddress[7]) );
  AOI22X1 U4613 ( .A(n4074), .B(instructionOrData), .C(n1034), .D(n4350), .Y(
        memoryAddress[8]) );
  AOI22X1 U4614 ( .A(n4072), .B(instructionOrData), .C(n1034), .D(n4351), .Y(
        memoryAddress[9]) );
  AOI22X1 U4615 ( .A(n4070), .B(instructionOrData), .C(n1034), .D(n4352), .Y(
        memoryAddress[10]) );
  AOI22X1 U4616 ( .A(n4068), .B(instructionOrData), .C(n1034), .D(n4353), .Y(
        memoryAddress[11]) );
  AOI22X1 U4617 ( .A(n4066), .B(instructionOrData), .C(n1034), .D(n4354), .Y(
        memoryAddress[12]) );
  AOI22X1 U4618 ( .A(n4064), .B(instructionOrData), .C(n1034), .D(n4355), .Y(
        memoryAddress[13]) );
  AOI22X1 U4619 ( .A(n4062), .B(instructionOrData), .C(n1034), .D(n4356), .Y(
        memoryAddress[14]) );
  AOI22X1 U4620 ( .A(n4060), .B(instructionOrData), .C(n1034), .D(n4357), .Y(
        memoryAddress[15]) );
  NOR3X1 U4621 ( .A(n3720), .B(n2222), .C(n2223), .Y(n4373) );
  OAI21X1 U4622 ( .A(n3724), .B(fpuReady), .C(n4366), .Y(n4374) );
  AOI21X1 U4623 ( .A(n61), .B(n4365), .C(n2212), .Y(n4375) );
endmodule

